magic
tech sky130A
magscale 1 2
timestamp 1649149387
<< obsli1 >>
rect 1104 2159 59064 59857
<< obsm1 >>
rect 14 1164 59970 59968
<< metal2 >>
rect 1306 61602 1362 62402
rect 3882 61602 3938 62402
rect 6458 61602 6514 62402
rect 9034 61602 9090 62402
rect 11610 61602 11666 62402
rect 13542 61602 13598 62402
rect 16118 61602 16174 62402
rect 18694 61602 18750 62402
rect 21270 61602 21326 62402
rect 23846 61602 23902 62402
rect 25778 61602 25834 62402
rect 28354 61602 28410 62402
rect 30930 61602 30986 62402
rect 33506 61602 33562 62402
rect 36082 61602 36138 62402
rect 38014 61602 38070 62402
rect 40590 61602 40646 62402
rect 43166 61602 43222 62402
rect 45742 61602 45798 62402
rect 48318 61602 48374 62402
rect 50250 61602 50306 62402
rect 52826 61602 52882 62402
rect 55402 61602 55458 62402
rect 57978 61602 58034 62402
rect 59910 61602 59966 62402
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 7102 0 7158 800
rect 9678 0 9734 800
rect 11610 0 11666 800
rect 14186 0 14242 800
rect 16762 0 16818 800
rect 19338 0 19394 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 26422 0 26478 800
rect 28998 0 29054 800
rect 31574 0 31630 800
rect 34150 0 34206 800
rect 36082 0 36138 800
rect 38658 0 38714 800
rect 41234 0 41290 800
rect 43810 0 43866 800
rect 46386 0 46442 800
rect 48318 0 48374 800
rect 50894 0 50950 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 58622 0 58678 800
<< obsm2 >>
rect 20 61546 1250 61985
rect 1418 61546 3826 61985
rect 3994 61546 6402 61985
rect 6570 61546 8978 61985
rect 9146 61546 11554 61985
rect 11722 61546 13486 61985
rect 13654 61546 16062 61985
rect 16230 61546 18638 61985
rect 18806 61546 21214 61985
rect 21382 61546 23790 61985
rect 23958 61546 25722 61985
rect 25890 61546 28298 61985
rect 28466 61546 30874 61985
rect 31042 61546 33450 61985
rect 33618 61546 36026 61985
rect 36194 61546 37958 61985
rect 38126 61546 40534 61985
rect 40702 61546 43110 61985
rect 43278 61546 45686 61985
rect 45854 61546 48262 61985
rect 48430 61546 50194 61985
rect 50362 61546 52770 61985
rect 52938 61546 55346 61985
rect 55514 61546 57922 61985
rect 58090 61546 59854 61985
rect 20 856 59964 61546
rect 130 31 1894 856
rect 2062 31 4470 856
rect 4638 31 7046 856
rect 7214 31 9622 856
rect 9790 31 11554 856
rect 11722 31 14130 856
rect 14298 31 16706 856
rect 16874 31 19282 856
rect 19450 31 21858 856
rect 22026 31 23790 856
rect 23958 31 26366 856
rect 26534 31 28942 856
rect 29110 31 31518 856
rect 31686 31 34094 856
rect 34262 31 36026 856
rect 36194 31 38602 856
rect 38770 31 41178 856
rect 41346 31 43754 856
rect 43922 31 46330 856
rect 46498 31 48262 856
rect 48430 31 50838 856
rect 51006 31 53414 856
rect 53582 31 55990 856
rect 56158 31 58566 856
rect 58734 31 59964 856
<< metal3 >>
rect 0 61888 800 62008
rect 59458 59848 60258 59968
rect 0 59168 800 59288
rect 59458 57128 60258 57248
rect 0 56448 800 56568
rect 59458 54408 60258 54528
rect 0 53728 800 53848
rect 59458 51688 60258 51808
rect 0 51008 800 51128
rect 59458 49648 60258 49768
rect 0 48968 800 49088
rect 59458 46928 60258 47048
rect 0 46248 800 46368
rect 59458 44208 60258 44328
rect 0 43528 800 43648
rect 59458 41488 60258 41608
rect 0 40808 800 40928
rect 59458 38768 60258 38888
rect 0 38088 800 38208
rect 59458 36728 60258 36848
rect 0 36048 800 36168
rect 59458 34008 60258 34128
rect 0 33328 800 33448
rect 59458 31288 60258 31408
rect 0 30608 800 30728
rect 59458 28568 60258 28688
rect 0 27888 800 28008
rect 59458 25848 60258 25968
rect 0 25168 800 25288
rect 59458 23808 60258 23928
rect 0 23128 800 23248
rect 59458 21088 60258 21208
rect 0 20408 800 20528
rect 59458 18368 60258 18488
rect 0 17688 800 17808
rect 59458 15648 60258 15768
rect 0 14968 800 15088
rect 59458 12928 60258 13048
rect 0 12248 800 12368
rect 59458 10888 60258 11008
rect 0 10208 800 10328
rect 59458 8168 60258 8288
rect 0 7488 800 7608
rect 59458 5448 60258 5568
rect 0 4768 800 4888
rect 59458 2728 60258 2848
rect 0 2048 800 2168
rect 59458 8 60258 128
<< obsm3 >>
rect 880 61808 59458 61981
rect 800 60048 59458 61808
rect 800 59768 59378 60048
rect 800 59368 59458 59768
rect 880 59088 59458 59368
rect 800 57328 59458 59088
rect 800 57048 59378 57328
rect 800 56648 59458 57048
rect 880 56368 59458 56648
rect 800 54608 59458 56368
rect 800 54328 59378 54608
rect 800 53928 59458 54328
rect 880 53648 59458 53928
rect 800 51888 59458 53648
rect 800 51608 59378 51888
rect 800 51208 59458 51608
rect 880 50928 59458 51208
rect 800 49848 59458 50928
rect 800 49568 59378 49848
rect 800 49168 59458 49568
rect 880 48888 59458 49168
rect 800 47128 59458 48888
rect 800 46848 59378 47128
rect 800 46448 59458 46848
rect 880 46168 59458 46448
rect 800 44408 59458 46168
rect 800 44128 59378 44408
rect 800 43728 59458 44128
rect 880 43448 59458 43728
rect 800 41688 59458 43448
rect 800 41408 59378 41688
rect 800 41008 59458 41408
rect 880 40728 59458 41008
rect 800 38968 59458 40728
rect 800 38688 59378 38968
rect 800 38288 59458 38688
rect 880 38008 59458 38288
rect 800 36928 59458 38008
rect 800 36648 59378 36928
rect 800 36248 59458 36648
rect 880 35968 59458 36248
rect 800 34208 59458 35968
rect 800 33928 59378 34208
rect 800 33528 59458 33928
rect 880 33248 59458 33528
rect 800 31488 59458 33248
rect 800 31208 59378 31488
rect 800 30808 59458 31208
rect 880 30528 59458 30808
rect 800 28768 59458 30528
rect 800 28488 59378 28768
rect 800 28088 59458 28488
rect 880 27808 59458 28088
rect 800 26048 59458 27808
rect 800 25768 59378 26048
rect 800 25368 59458 25768
rect 880 25088 59458 25368
rect 800 24008 59458 25088
rect 800 23728 59378 24008
rect 800 23328 59458 23728
rect 880 23048 59458 23328
rect 800 21288 59458 23048
rect 800 21008 59378 21288
rect 800 20608 59458 21008
rect 880 20328 59458 20608
rect 800 18568 59458 20328
rect 800 18288 59378 18568
rect 800 17888 59458 18288
rect 880 17608 59458 17888
rect 800 15848 59458 17608
rect 800 15568 59378 15848
rect 800 15168 59458 15568
rect 880 14888 59458 15168
rect 800 13128 59458 14888
rect 800 12848 59378 13128
rect 800 12448 59458 12848
rect 880 12168 59458 12448
rect 800 11088 59458 12168
rect 800 10808 59378 11088
rect 800 10408 59458 10808
rect 880 10128 59458 10408
rect 800 8368 59458 10128
rect 800 8088 59378 8368
rect 800 7688 59458 8088
rect 880 7408 59458 7688
rect 800 5648 59458 7408
rect 800 5368 59378 5648
rect 800 4968 59458 5368
rect 880 4688 59458 4968
rect 800 2928 59458 4688
rect 800 2648 59378 2928
rect 800 2248 59458 2648
rect 880 1968 59458 2248
rect 800 208 59458 1968
rect 800 35 59378 208
<< metal4 >>
rect 4208 2128 4528 59888
rect 19568 2128 19888 59888
rect 34928 2128 35248 59888
rect 50288 2128 50608 59888
<< obsm4 >>
rect 1899 2211 4128 58037
rect 4608 2211 19488 58037
rect 19968 2211 34848 58037
rect 35328 2211 50208 58037
rect 50688 2211 55141 58037
<< metal5 >>
rect 1104 51252 59064 51572
rect 1104 35934 59064 36254
rect 1104 20616 59064 20936
rect 1104 5298 59064 5618
<< obsm5 >>
rect 15020 6980 31164 10700
<< labels >>
rlabel metal2 s 7102 0 7158 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 40590 61602 40646 62402 6 A[10]
port 2 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 A[11]
port 3 nsew signal input
rlabel metal2 s 57978 61602 58034 62402 6 A[12]
port 4 nsew signal input
rlabel metal3 s 59458 51688 60258 51808 6 A[13]
port 5 nsew signal input
rlabel metal3 s 59458 38768 60258 38888 6 A[14]
port 6 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 A[15]
port 7 nsew signal input
rlabel metal2 s 21270 61602 21326 62402 6 A[16]
port 8 nsew signal input
rlabel metal2 s 23846 61602 23902 62402 6 A[17]
port 9 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 A[18]
port 10 nsew signal input
rlabel metal3 s 59458 59848 60258 59968 6 A[19]
port 11 nsew signal input
rlabel metal3 s 59458 15648 60258 15768 6 A[1]
port 12 nsew signal input
rlabel metal3 s 59458 49648 60258 49768 6 A[20]
port 13 nsew signal input
rlabel metal2 s 18694 61602 18750 62402 6 A[21]
port 14 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 A[22]
port 15 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 A[23]
port 16 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 A[24]
port 17 nsew signal input
rlabel metal3 s 59458 57128 60258 57248 6 A[25]
port 18 nsew signal input
rlabel metal2 s 16118 61602 16174 62402 6 A[26]
port 19 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 A[27]
port 20 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 A[28]
port 21 nsew signal input
rlabel metal3 s 59458 23808 60258 23928 6 A[29]
port 22 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 A[2]
port 23 nsew signal input
rlabel metal3 s 59458 34008 60258 34128 6 A[30]
port 24 nsew signal input
rlabel metal3 s 59458 18368 60258 18488 6 A[31]
port 25 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 A[3]
port 26 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 A[4]
port 27 nsew signal input
rlabel metal3 s 59458 46928 60258 47048 6 A[5]
port 28 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 A[6]
port 29 nsew signal input
rlabel metal3 s 59458 8168 60258 8288 6 A[7]
port 30 nsew signal input
rlabel metal3 s 59458 54408 60258 54528 6 A[8]
port 31 nsew signal input
rlabel metal2 s 38014 61602 38070 62402 6 A[9]
port 32 nsew signal input
rlabel metal2 s 28354 61602 28410 62402 6 B[0]
port 33 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 B[10]
port 34 nsew signal input
rlabel metal2 s 50250 61602 50306 62402 6 B[11]
port 35 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 B[12]
port 36 nsew signal input
rlabel metal3 s 59458 8 60258 128 6 B[13]
port 37 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 B[14]
port 38 nsew signal input
rlabel metal2 s 25778 61602 25834 62402 6 B[15]
port 39 nsew signal input
rlabel metal2 s 33506 61602 33562 62402 6 B[16]
port 40 nsew signal input
rlabel metal2 s 52826 61602 52882 62402 6 B[17]
port 41 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 B[18]
port 42 nsew signal input
rlabel metal3 s 59458 44208 60258 44328 6 B[19]
port 43 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 B[1]
port 44 nsew signal input
rlabel metal2 s 36082 61602 36138 62402 6 B[20]
port 45 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 B[21]
port 46 nsew signal input
rlabel metal3 s 59458 10888 60258 11008 6 B[22]
port 47 nsew signal input
rlabel metal3 s 59458 31288 60258 31408 6 B[23]
port 48 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 B[24]
port 49 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 B[25]
port 50 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 B[26]
port 51 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 B[27]
port 52 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 B[28]
port 53 nsew signal input
rlabel metal2 s 6458 61602 6514 62402 6 B[29]
port 54 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 B[2]
port 55 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 B[30]
port 56 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 B[31]
port 57 nsew signal input
rlabel metal3 s 59458 25848 60258 25968 6 B[3]
port 58 nsew signal input
rlabel metal3 s 59458 12928 60258 13048 6 B[4]
port 59 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 B[5]
port 60 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 B[6]
port 61 nsew signal input
rlabel metal3 s 59458 2728 60258 2848 6 B[7]
port 62 nsew signal input
rlabel metal2 s 9034 61602 9090 62402 6 B[8]
port 63 nsew signal input
rlabel metal3 s 59458 21088 60258 21208 6 B[9]
port 64 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 F[0]
port 65 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 F[10]
port 66 nsew signal output
rlabel metal3 s 59458 41488 60258 41608 6 F[11]
port 67 nsew signal output
rlabel metal2 s 11610 61602 11666 62402 6 F[12]
port 68 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 F[13]
port 69 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 F[14]
port 70 nsew signal output
rlabel metal2 s 18 0 74 800 6 F[15]
port 71 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 F[16]
port 72 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 F[17]
port 73 nsew signal output
rlabel metal2 s 30930 61602 30986 62402 6 F[18]
port 74 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 F[19]
port 75 nsew signal output
rlabel metal2 s 1306 61602 1362 62402 6 F[1]
port 76 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 F[20]
port 77 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 F[21]
port 78 nsew signal output
rlabel metal2 s 55402 61602 55458 62402 6 F[22]
port 79 nsew signal output
rlabel metal2 s 43166 61602 43222 62402 6 F[23]
port 80 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 F[24]
port 81 nsew signal output
rlabel metal2 s 59910 61602 59966 62402 6 F[25]
port 82 nsew signal output
rlabel metal3 s 59458 5448 60258 5568 6 F[26]
port 83 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 F[27]
port 84 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 F[28]
port 85 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 F[29]
port 86 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 F[2]
port 87 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 F[30]
port 88 nsew signal output
rlabel metal3 s 59458 36728 60258 36848 6 F[31]
port 89 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 F[3]
port 90 nsew signal output
rlabel metal2 s 48318 61602 48374 62402 6 F[4]
port 91 nsew signal output
rlabel metal2 s 45742 61602 45798 62402 6 F[5]
port 92 nsew signal output
rlabel metal2 s 3882 61602 3938 62402 6 F[6]
port 93 nsew signal output
rlabel metal2 s 13542 61602 13598 62402 6 F[7]
port 94 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 F[8]
port 95 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 F[9]
port 96 nsew signal output
rlabel metal5 s 1104 20616 59064 20936 6 VGND
port 97 nsew ground input
rlabel metal5 s 1104 51252 59064 51572 6 VGND
port 97 nsew ground input
rlabel metal4 s 19568 2128 19888 59888 6 VGND
port 97 nsew ground input
rlabel metal4 s 50288 2128 50608 59888 6 VGND
port 97 nsew ground input
rlabel metal5 s 1104 5298 59064 5618 6 VPWR
port 98 nsew power input
rlabel metal5 s 1104 35934 59064 36254 6 VPWR
port 98 nsew power input
rlabel metal4 s 4208 2128 4528 59888 6 VPWR
port 98 nsew power input
rlabel metal4 s 34928 2128 35248 59888 6 VPWR
port 98 nsew power input
rlabel metal3 s 0 53728 800 53848 6 clk
port 99 nsew signal input
rlabel metal3 s 59458 28568 60258 28688 6 rst
port 100 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60258 62402
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14178468
string GDS_FILE /openlane/designs/MULTI_32bit/runs/RUN_2022.04.05_08.50.19/results/finishing/MULTI_32bit.magic.gds
string GDS_START 985846
<< end >>

