
.SUBCKT sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Y C2 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 net62 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net62 C2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net36 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net36 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net31 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net35 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net31 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Y A net35 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
rI12 VGND LO short
rI11 HI VPWR short
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net118 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net118 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net181 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net181 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net83 net121 net109 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net109 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net102 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net94 M1 net102 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net121 clkneg net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net83 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net82 net83 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net121 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net166 net83 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net83 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net121 clkpos net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net83 net121 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net145 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net145 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net145 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net83 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net121 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net129 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net80 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net129 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net97 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net89 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net89 S1 net97 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net80 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net141 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net141 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net192 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net192 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net156 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net141 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net141 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net128 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net111 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net96 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net88 S1 net96 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net111 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net140 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net140 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net191 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net191 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net168 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net168 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net155 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net140 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net140 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=1 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=5 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=5 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net121 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net121 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net112 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net56 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net112 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net56 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net52 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net52 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net112 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net112 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net107 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net107 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net87 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net87 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net53 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net53 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net44 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net96 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net76 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net76 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net55 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net55 net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 X net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net55 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net55 net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 X net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
MMIN1 Ab X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 net43 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net43 net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 X net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 net43 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net43 net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net56 net48 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net52 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net48 net44 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net44 net52 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net56 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net56 net48 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net48 net44 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net44 net52 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net52 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
MI14 net124 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net124 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net68 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net92 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net92 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net85 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net85 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net68 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Q_N S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net193 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net193 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net148 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net168 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net168 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net161 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net161 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net148 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net141 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net141 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Q_N S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
MI14 net115 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net115 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net59 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net79 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net83 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net83 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net79 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net76 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net76 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net59 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net175 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net175 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net172 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net148 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net148 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net172 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net128 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj31 sndNCINn3 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND A sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR A sndPCINp3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 sndPCINp3 CIN majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj31 sndPCINp3 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
MMIN2 COUT net195 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net123 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb mid2 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Bb mid1 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb mid2 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb mid1 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 CIbb CIb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 CIb CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Ab2 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 Abb2 Ab2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 Ab1 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb2 B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab1 Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb2 Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab1 B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT net195 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM net123 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb mid1 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb mid2 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb mid1 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb mid2 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 CIbb CIb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 CIb CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 Ab2 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 Abb2 Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 Ab1 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb2 Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab1 B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb2 B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab1 Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMIP3 SUM net144 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bbb Bb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CINb1 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CINbb2 CINb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CINb2 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CINbb2 mid2 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CINb2 mid1 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bbb mid2 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CINb1 mid1 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net144 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CINb1 mid2 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CINb1 CIN VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CINbb2 CINb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CINb2 CIN VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CINbb2 mid1 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CINb2 mid2 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bbb mid1 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bbb Bb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
MMIP3 SUM net146 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bb2 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb1 mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb1 mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CIb1 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CIbb2 CIb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CIb2 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb1 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb2 mid2 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb2 mid1 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb2 mid2 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb1 mid1 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net146 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb1 mid2 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb1 mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb1 mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CIb1 CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CIbb2 CIb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CIb2 CI VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb1 B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb2 mid1 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb2 mid2 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bb2 mid1 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bb2 B VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
MI2 net29 SHORT net25 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net25 SHORT net24 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VPWR SHORT net29 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net24 SHORT net16 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net16 SHORT VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net36 A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 sndA SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 net36 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
MI8 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net36 sleepb VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 sleepb SLEEP VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 sleepb sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 sleepb SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 sndA A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
MI23 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 VPWR net44 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 net56 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA net56 net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 net56 SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net44 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X net44 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net44 net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA A net36 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 VPWR net36 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net36 SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
MI677 Q s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 sleepneg sleeppos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI674 net39 s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 s0 sleepneg net49 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net49 D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 sleeppos net38 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net38 net39 VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 sleeppos SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 sleeppos SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 sleepneg sleeppos VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
MI662 net86 net39 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 sleepneg net86 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net39 s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 s0 sleeppos net69 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net69 D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA net58 net66 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net58 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab net66 KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net66 SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 net66 net58 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net58 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Ab net66 VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
MI2 net72 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 cross1 net72 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Ab A LOWLVPWR LOWLVPWR pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 X net60 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 net60 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 cross1 Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net72 A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 X net60 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 net60 cross1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
XI1 net59 LO VGND VNB VPB VPWR / sky130_fd_sc_hd__conb_1
XI6 nor2right invright VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI7 nor2left invleft VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI4 nd2right nd2right nor2right VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI5 nd2left nd2left nor2left VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI2 LO LO nd2right VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
XI3 LO LO nd2left VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.7 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net29 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net29 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net29 X short
.ENDS




.SUBCKT sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net33 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net33 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net33 X short
rI120 VGND met5vgnd short
rI119 VPWR met5vpwr short
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net153 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net153 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net128 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net103 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net103 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net87 net153 net117 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net117 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net110 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net98 M1 net110 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net153 clkneg net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net87 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net93 net87 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net153 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net87 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net87 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net153 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net87 net153 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net87 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net153 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net83 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net83 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net159 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net159 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net138 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net199 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net199 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net98 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net98 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI27 net243 S1 net215 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net230 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net227 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net199 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net215 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net199 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net227 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net230 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net243 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net195 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net195 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net130 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net130 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net107 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI34 S0 clkpos net219 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net239 S1 net187 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net230 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net199 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net230 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net219 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net239 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net199 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net195 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net187 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net195 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net212 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net196 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net212 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net196 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net104 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net104 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net177 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net160 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net177 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net160 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net196 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net189 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net196 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net189 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net138 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net123 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net123 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net235 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net235 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net203 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net203 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net240 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net240 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net180 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net180 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net103 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net103 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net179 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net179 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net135 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net135 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net227 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net227 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net190 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net190 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net163 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net163 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS

















































































































































.subckt MULTI_32bit A[0] A[10] A[11] A[12] A[13] A[14] A[15] A[16] A[17] A[18] A[19]
+ A[1] A[20] A[21] A[22] A[23] A[24] A[25] A[26] A[27] A[28] A[29] A[2] A[30] A[31]
+ A[3] A[4] A[5] A[6] A[7] A[8] A[9] B[0] B[10] B[11] B[12] B[13] B[14] B[15] B[16]
+ B[17] B[18] B[19] B[1] B[20] B[21] B[22] B[23] B[24] B[25] B[26] B[27] B[28] B[29]
+ B[2] B[30] B[31] B[3] B[4] B[5] B[6] B[7] B[8] B[9] F[0] F[10] F[11] F[12] F[13]
+ F[14] F[15] F[16] F[17] F[18] F[19] F[1] F[20] F[21] F[22] F[23] F[24] F[25] F[26]
+ F[27] F[28] F[29] F[2] F[30] F[31] F[3] F[4] F[5] F[6] F[7] F[8] F[9] VGND VPWR
+ clk rst
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7963_ _7963_/A _7963_/B VGND VGND VPWR VPWR _7974_/A sky130_fd_sc_hd__xnor2_1
X_6914_ _7029_/B VGND VGND VPWR VPWR _6914_/Y sky130_fd_sc_hd__inv_2
X_7894_ _7894_/A _7894_/B VGND VGND VPWR VPWR _7897_/A sky130_fd_sc_hd__xnor2_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6845_ _6845_/A _6845_/B _6845_/C VGND VGND VPWR VPWR _6845_/X sky130_fd_sc_hd__and3_1
X_6776_ _9179_/Q VGND VGND VPWR VPWR _7119_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_8515_ _8337_/A _8351_/B _8516_/B _8587_/A VGND VGND VPWR VPWR _8518_/A sky130_fd_sc_hd__a22oi_1
XFILLER_10_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5727_ _4780_/A _5726_/X _5727_/S VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__mux2_1
X_8446_ _8447_/A _8447_/B _8447_/C VGND VGND VPWR VPWR _8556_/A sky130_fd_sc_hd__o21a_1
X_5658_ _4846_/A _5119_/A _5656_/Y _5657_/X _5140_/A VGND VGND VPWR VPWR _5658_/X
+ sky130_fd_sc_hd__a221o_1
X_8377_ _8377_/A _8377_/B VGND VGND VPWR VPWR _8397_/A sky130_fd_sc_hd__xor2_1
X_5589_ _5249_/A _5389_/A _5258_/A VGND VGND VPWR VPWR _5589_/Y sky130_fd_sc_hd__a21oi_1
X_4609_ _9104_/Q VGND VGND VPWR VPWR _5735_/S sky130_fd_sc_hd__inv_2
XFILLER_89_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7328_ _7328_/A _7328_/B VGND VGND VPWR VPWR _7329_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7259_ _7259_/A _7259_/B _9180_/Q _7259_/D VGND VGND VPWR VPWR _7260_/B sky130_fd_sc_hd__and4_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4960_ _4960_/A _4960_/B _4963_/B VGND VGND VPWR VPWR _4960_/X sky130_fd_sc_hd__and3_1
XFILLER_83_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4891_ _4891_/A VGND VGND VPWR VPWR _4891_/X sky130_fd_sc_hd__clkbuf_2
X_6630_ _8519_/A VGND VGND VPWR VPWR _8584_/A sky130_fd_sc_hd__buf_4
X_6561_ _6558_/X _6649_/B _6478_/B _6480_/X VGND VGND VPWR VPWR _6562_/B sky130_fd_sc_hd__o211a_1
X_8300_ _8393_/B _8300_/B VGND VGND VPWR VPWR _8304_/A sky130_fd_sc_hd__or2_1
X_5512_ _4849_/A _5179_/A _4846_/A VGND VGND VPWR VPWR _5512_/Y sky130_fd_sc_hd__a21oi_1
X_6492_ _7148_/D VGND VGND VPWR VPWR _7604_/D sky130_fd_sc_hd__clkbuf_2
X_8231_ _8231_/A _8231_/B VGND VGND VPWR VPWR _8232_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5443_ _5382_/X _5278_/X _5414_/X VGND VGND VPWR VPWR _5443_/Y sky130_fd_sc_hd__a21oi_1
X_8162_ _8162_/A _8162_/B VGND VGND VPWR VPWR _8164_/B sky130_fd_sc_hd__xnor2_1
X_5374_ _5142_/X _5248_/Y _5154_/X VGND VGND VPWR VPWR _5374_/Y sky130_fd_sc_hd__a21oi_1
X_7113_ _9182_/Q VGND VGND VPWR VPWR _7640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8093_ _8093_/A _8150_/D VGND VGND VPWR VPWR _8094_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7044_ _7044_/A _7044_/B VGND VGND VPWR VPWR _7143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8995_ _8993_/X _9018_/A _8948_/A _8952_/B VGND VGND VPWR VPWR _8995_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7946_ _7946_/A _7946_/B _7945_/X VGND VGND VPWR VPWR _7948_/A sky130_fd_sc_hd__or3b_1
XFILLER_55_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7877_ _7877_/A _7976_/A VGND VGND VPWR VPWR _7957_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6828_ _6828_/A _7824_/B VGND VGND VPWR VPWR _6829_/B sky130_fd_sc_hd__nand2_2
X_6759_ _7148_/A _7040_/A _6759_/C _6927_/D VGND VGND VPWR VPWR _6762_/A sky130_fd_sc_hd__and4_1
XFILLER_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8429_ _8510_/A _8429_/B VGND VGND VPWR VPWR _8430_/B sky130_fd_sc_hd__and2b_1
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5090_ _4940_/C _4998_/A _5040_/A _5740_/S VGND VGND VPWR VPWR _5090_/X sky130_fd_sc_hd__a31o_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8780_ _8780_/A _8780_/B _8887_/A VGND VGND VPWR VPWR _8836_/A sky130_fd_sc_hd__and3_1
X_7800_ _7699_/A _7699_/B _7703_/B VGND VGND VPWR VPWR _7800_/Y sky130_fd_sc_hd__a21oi_1
X_5992_ _5979_/A _5979_/B _5979_/C VGND VGND VPWR VPWR _6037_/C sky130_fd_sc_hd__a21o_1
XFILLER_91_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7731_ _7731_/A _7731_/B VGND VGND VPWR VPWR _7739_/A sky130_fd_sc_hd__xnor2_2
X_4943_ _4943_/A _4943_/B VGND VGND VPWR VPWR _5093_/A sky130_fd_sc_hd__and2_2
X_7662_ _7661_/A _7661_/B _7660_/Y VGND VGND VPWR VPWR _7784_/A sky130_fd_sc_hd__o21ba_2
XFILLER_60_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6613_ _6614_/B _6691_/A _6614_/A VGND VGND VPWR VPWR _6615_/A sky130_fd_sc_hd__a21o_1
X_4874_ _4872_/X _4873_/Y _4874_/S VGND VGND VPWR VPWR _4874_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7593_ _7594_/A _7594_/B VGND VGND VPWR VPWR _7593_/X sky130_fd_sc_hd__and2_1
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _9212_/CLK sky130_fd_sc_hd__clkbuf_2
X_6544_ _6543_/B _6616_/A _6543_/A VGND VGND VPWR VPWR _6545_/B sky130_fd_sc_hd__a21o_1
X_6475_ _6560_/B _6475_/B VGND VGND VPWR VPWR _6476_/C sky130_fd_sc_hd__xnor2_1
X_8214_ _8898_/B VGND VGND VPWR VPWR _8933_/B sky130_fd_sc_hd__buf_2
X_5426_ _5287_/X _5187_/X _5422_/X _5425_/Y VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__a22o_1
X_9194_ _9219_/CLK _9194_/D VGND VGND VPWR VPWR _9194_/Q sky130_fd_sc_hd__dfxtp_4
X_8145_ _8254_/A _8145_/B VGND VGND VPWR VPWR _8168_/A sky130_fd_sc_hd__and2_1
X_5357_ _5245_/X _5356_/X _5427_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8076_ _8076_/A _8076_/B VGND VGND VPWR VPWR _8078_/C sky130_fd_sc_hd__xnor2_1
X_5288_ _5362_/A _5559_/B VGND VGND VPWR VPWR _5288_/X sky130_fd_sc_hd__or2_1
XFILLER_87_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7027_ _7027_/A _7027_/B _7141_/A VGND VGND VPWR VPWR _7141_/B sky130_fd_sc_hd__nand3_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8978_ _8978_/A _8978_/B _9002_/A VGND VGND VPWR VPWR _8979_/A sky130_fd_sc_hd__and3_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7929_ _7929_/A _7929_/B VGND VGND VPWR VPWR _7932_/A sky130_fd_sc_hd__xor2_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4590_ _4839_/A VGND VGND VPWR VPWR _4591_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR clkbuf_4_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6260_ _6260_/A _6351_/B VGND VGND VPWR VPWR _6352_/B sky130_fd_sc_hd__xnor2_1
X_6191_ _6361_/D VGND VGND VPWR VPWR _8091_/B sky130_fd_sc_hd__clkbuf_2
X_5211_ _5211_/A VGND VGND VPWR VPWR _5212_/A sky130_fd_sc_hd__inv_2
X_5142_ _5151_/A VGND VGND VPWR VPWR _5142_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5073_ _5074_/A _5080_/C _5074_/B VGND VGND VPWR VPWR _5073_/Y sky130_fd_sc_hd__o21ai_1
X_8901_ _8901_/A _8945_/B VGND VGND VPWR VPWR _8902_/B sky130_fd_sc_hd__nand2_1
X_8832_ _8832_/A _8832_/B VGND VGND VPWR VPWR _8937_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8763_ _8763_/A _8825_/A VGND VGND VPWR VPWR _8776_/A sky130_fd_sc_hd__and2_1
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5975_ _5968_/A _5968_/B _5968_/C VGND VGND VPWR VPWR _5976_/C sky130_fd_sc_hd__a21o_1
XFILLER_40_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8694_ _8694_/A _8750_/A _8694_/C VGND VGND VPWR VPWR _8761_/A sky130_fd_sc_hd__and3_1
X_7714_ _7588_/A _7714_/B VGND VGND VPWR VPWR _7714_/X sky130_fd_sc_hd__and2b_1
XFILLER_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4926_ _4925_/A _4950_/B _5730_/S VGND VGND VPWR VPWR _4926_/X sky130_fd_sc_hd__a21o_1
X_7645_ _7645_/A _7769_/A _7645_/C VGND VGND VPWR VPWR _7651_/B sky130_fd_sc_hd__and3_1
XFILLER_20_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4857_ _4857_/A VGND VGND VPWR VPWR _5007_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7576_ _7576_/A _7576_/B VGND VGND VPWR VPWR _7577_/B sky130_fd_sc_hd__and2_1
X_6527_ _9176_/Q VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4788_ _5621_/A _4786_/X _4787_/Y _5222_/A VGND VGND VPWR VPWR _4788_/X sky130_fd_sc_hd__a211o_1
X_6458_ _6458_/A _6458_/B _6458_/C VGND VGND VPWR VPWR _6512_/B sky130_fd_sc_hd__nand3_1
X_6389_ _7222_/C VGND VGND VPWR VPWR _7604_/C sky130_fd_sc_hd__clkbuf_2
X_5409_ _5249_/X _5179_/X _5258_/X VGND VGND VPWR VPWR _5409_/Y sky130_fd_sc_hd__a21oi_1
X_9177_ _9220_/CLK input7/X VGND VGND VPWR VPWR _9177_/Q sky130_fd_sc_hd__dfxtp_4
X_8128_ _8128_/A _8128_/B VGND VGND VPWR VPWR _8128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8059_ _8058_/A _8058_/B _8057_/X VGND VGND VPWR VPWR _8060_/B sky130_fd_sc_hd__o21bai_2
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5760_ _5632_/X _4889_/X _5759_/X _5698_/S VGND VGND VPWR VPWR _5760_/X sky130_fd_sc_hd__o31a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5691_ _5136_/X _5690_/X _5691_/S VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__mux2_1
X_4711_ _4693_/Y _4709_/X _5728_/S VGND VGND VPWR VPWR _4711_/X sky130_fd_sc_hd__mux2_1
X_7430_ _7696_/C VGND VGND VPWR VPWR _7918_/A sky130_fd_sc_hd__clkbuf_2
X_4642_ _4642_/A VGND VGND VPWR VPWR _4643_/A sky130_fd_sc_hd__clkbuf_2
X_7361_ _7358_/Y _7482_/A _7361_/C _7756_/A VGND VGND VPWR VPWR _7482_/B sky130_fd_sc_hd__and4bb_1
X_4573_ _4573_/A VGND VGND VPWR VPWR _4573_/X sky130_fd_sc_hd__clkbuf_2
X_6312_ _7129_/B VGND VGND VPWR VPWR _7604_/B sky130_fd_sc_hd__clkbuf_2
X_9100_ _9221_/CLK _9100_/D VGND VGND VPWR VPWR _9100_/Q sky130_fd_sc_hd__dfxtp_1
X_7292_ _7295_/D VGND VGND VPWR VPWR _7292_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9031_ _9031_/A _9031_/B VGND VGND VPWR VPWR _9032_/B sky130_fd_sc_hd__nor2_1
X_6243_ _6335_/A _6335_/B VGND VGND VPWR VPWR _6245_/A sky130_fd_sc_hd__xor2_1
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6174_ _7293_/B _6907_/A _7986_/A _6251_/A VGND VGND VPWR VPWR _6175_/B sky130_fd_sc_hd__a22oi_2
XFILLER_97_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5125_ _5125_/A VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5056_ _4845_/A _5052_/A _5067_/A _5053_/A VGND VGND VPWR VPWR _5056_/X sky130_fd_sc_hd__a31o_1
X_8815_ _8813_/X _8815_/B VGND VGND VPWR VPWR _8817_/A sky130_fd_sc_hd__and2b_1
X_8746_ _8746_/A _8806_/B _8746_/C VGND VGND VPWR VPWR _8814_/A sky130_fd_sc_hd__and3_1
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5958_ _5958_/A VGND VGND VPWR VPWR _9073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4909_ _4937_/B VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__clkbuf_2
X_8677_ _8677_/A _8733_/A _8842_/A _8733_/D VGND VGND VPWR VPWR _8678_/B sky130_fd_sc_hd__and4_1
X_5889_ _6825_/B VGND VGND VPWR VPWR _6359_/A sky130_fd_sc_hd__clkbuf_2
X_7628_ _7628_/A _8091_/C VGND VGND VPWR VPWR _7629_/B sky130_fd_sc_hd__nand2_1
X_7559_ _7559_/A _7559_/B _7558_/Y VGND VGND VPWR VPWR _7561_/A sky130_fd_sc_hd__nor3b_1
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_5 _9199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6930_ _6930_/A _6930_/B VGND VGND VPWR VPWR _7031_/B sky130_fd_sc_hd__xnor2_2
XFILLER_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6861_ _6861_/A _6861_/B VGND VGND VPWR VPWR _6862_/B sky130_fd_sc_hd__nor2_1
X_8600_ _8600_/A _8600_/B VGND VGND VPWR VPWR _8603_/A sky130_fd_sc_hd__xor2_1
X_6792_ _6671_/A _6670_/B _6670_/A VGND VGND VPWR VPWR _6883_/A sky130_fd_sc_hd__o21ba_1
XFILLER_50_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5812_ _5812_/A _5812_/B VGND VGND VPWR VPWR _5834_/A sky130_fd_sc_hd__xor2_4
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8531_ _8700_/A _8846_/B _8529_/Y _8530_/X VGND VGND VPWR VPWR _8533_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5743_ _5765_/B _5742_/X _5743_/S VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__mux2_1
X_8462_ _8756_/A _8832_/A _8390_/A _8387_/B VGND VGND VPWR VPWR _8473_/A sky130_fd_sc_hd__a31o_1
X_5674_ _5606_/X _5673_/X _5674_/S VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__mux2_1
X_8393_ _8393_/A _8393_/B _8392_/Y VGND VGND VPWR VPWR _8395_/A sky130_fd_sc_hd__or3b_1
X_4625_ _5765_/B _4621_/X _5282_/S VGND VGND VPWR VPWR _4625_/X sky130_fd_sc_hd__o21a_1
X_7413_ _7804_/B VGND VGND VPWR VPWR _8867_/B sky130_fd_sc_hd__clkbuf_4
X_7344_ _7342_/X _7234_/B _7340_/X _7341_/Y VGND VGND VPWR VPWR _7416_/A sky130_fd_sc_hd__a211oi_2
X_4556_ _4556_/A VGND VGND VPWR VPWR _5378_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7275_ _7274_/A _7274_/B _7274_/C VGND VGND VPWR VPWR _7277_/D sky130_fd_sc_hd__a21oi_4
XFILLER_103_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9014_ _9014_/A _9035_/A VGND VGND VPWR VPWR _9017_/A sky130_fd_sc_hd__and2_1
X_6226_ _7152_/B VGND VGND VPWR VPWR _7822_/A sky130_fd_sc_hd__clkbuf_2
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6157_/A _6157_/B VGND VGND VPWR VPWR _6161_/A sky130_fd_sc_hd__nor2_2
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _4687_/X _5107_/X _5098_/X VGND VGND VPWR VPWR _5108_/X sky130_fd_sc_hd__o21a_1
X_6088_ _6018_/A _6018_/B _6018_/C VGND VGND VPWR VPWR _6090_/C sky130_fd_sc_hd__a21bo_1
XFILLER_72_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5039_ _5080_/B VGND VGND VPWR VPWR _5040_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8729_ _8729_/A _8729_/B VGND VGND VPWR VPWR _8805_/A sky130_fd_sc_hd__or2_1
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput75 _9148_/Q VGND VGND VPWR VPWR F[19] sky130_fd_sc_hd__buf_2
Xoutput86 _9158_/Q VGND VGND VPWR VPWR F[29] sky130_fd_sc_hd__buf_2
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5390_ _5271_/X _5389_/X _4629_/A VGND VGND VPWR VPWR _5390_/Y sky130_fd_sc_hd__a21oi_1
X_7060_ _7073_/B _7060_/B VGND VGND VPWR VPWR _7061_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6011_ _6169_/A _7253_/B _9170_/Q _6240_/A VGND VGND VPWR VPWR _6013_/A sky130_fd_sc_hd__a22oi_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7962_ _8379_/A _7962_/B VGND VGND VPWR VPWR _7963_/B sky130_fd_sc_hd__nand2_1
X_6913_ _6913_/A _6913_/B _7029_/A VGND VGND VPWR VPWR _7029_/B sky130_fd_sc_hd__nand3_2
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7893_ _7893_/A _7893_/B VGND VGND VPWR VPWR _7894_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6844_ _6844_/A _6844_/B VGND VGND VPWR VPWR _6847_/A sky130_fd_sc_hd__or2_1
X_6775_ _6775_/A _7604_/B VGND VGND VPWR VPWR _6781_/A sky130_fd_sc_hd__nand2_1
X_8514_ _8514_/A _8435_/B VGND VGND VPWR VPWR _8525_/A sky130_fd_sc_hd__or2b_1
X_5726_ _4776_/A _4582_/A _5725_/X VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__a21o_1
X_8445_ _8445_/A _8525_/B VGND VGND VPWR VPWR _8447_/C sky130_fd_sc_hd__and2_1
X_5657_ _5252_/A _9087_/Q _4658_/A _9085_/Q _4706_/S VGND VGND VPWR VPWR _5657_/X
+ sky130_fd_sc_hd__o221a_1
X_8376_ _8498_/A _8850_/B VGND VGND VPWR VPWR _8377_/B sky130_fd_sc_hd__nand2_1
X_5588_ _4862_/X _5205_/A _5587_/X _4841_/A VGND VGND VPWR VPWR _5588_/X sky130_fd_sc_hd__a211o_1
X_4608_ _4637_/A _4608_/B VGND VGND VPWR VPWR _4608_/X sky130_fd_sc_hd__or2_1
X_7327_ _7327_/A _7327_/B _7327_/C _9206_/Q VGND VGND VPWR VPWR _7328_/B sky130_fd_sc_hd__and4_1
XFILLER_2_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4539_ _9107_/Q VGND VGND VPWR VPWR _5391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7258_ _7259_/A _7119_/D _7259_/D _7119_/B VGND VGND VPWR VPWR _7260_/A sky130_fd_sc_hd__a22oi_1
XFILLER_104_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6209_ _6210_/A _6210_/B _6210_/C VGND VGND VPWR VPWR _6211_/A sky130_fd_sc_hd__a21oi_1
X_7189_ _7187_/X _7571_/A _7189_/C _7189_/D VGND VGND VPWR VPWR _7190_/B sky130_fd_sc_hd__and4b_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4890_ _4889_/X _4873_/A _4538_/A VGND VGND VPWR VPWR _4890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6560_ _6560_/A _6560_/B _6560_/C VGND VGND VPWR VPWR _6649_/B sky130_fd_sc_hd__nor3_1
X_5511_ _5511_/A VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__clkbuf_2
X_6491_ _7327_/C VGND VGND VPWR VPWR _6493_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8230_ _8230_/A _8333_/A VGND VGND VPWR VPWR _8232_/A sky130_fd_sc_hd__nor2_1
X_5442_ _5367_/X _5208_/X _5440_/X _5441_/Y _5380_/X VGND VGND VPWR VPWR _5442_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8161_ _8236_/B _8161_/B VGND VGND VPWR VPWR _8162_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5373_ _5149_/X _5507_/A _5370_/Y _5372_/X _5151_/X VGND VGND VPWR VPWR _5373_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8092_ _8092_/A _8092_/B VGND VGND VPWR VPWR _8094_/A sky130_fd_sc_hd__nor2_1
X_7112_ _7253_/A _9178_/Q _7767_/C VGND VGND VPWR VPWR _7246_/A sky130_fd_sc_hd__and3_1
XFILLER_101_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7043_ _7043_/A _7043_/B VGND VGND VPWR VPWR _7044_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8994_ _8955_/A _9013_/A _8994_/C VGND VGND VPWR VPWR _9018_/A sky130_fd_sc_hd__and3b_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7945_ _8058_/B _7945_/B VGND VGND VPWR VPWR _7945_/X sky130_fd_sc_hd__or2_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7876_ _7876_/A _7876_/B VGND VGND VPWR VPWR _7976_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6827_ _9210_/Q VGND VGND VPWR VPWR _7824_/B sky130_fd_sc_hd__buf_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6758_ _7694_/A _7608_/A VGND VGND VPWR VPWR _6763_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6689_ _6689_/A _6689_/B _6810_/A VGND VGND VPWR VPWR _6810_/B sky130_fd_sc_hd__nand3_2
X_5709_ _4635_/A _5378_/X _5707_/X _5708_/Y _4607_/A VGND VGND VPWR VPWR _5709_/X
+ sky130_fd_sc_hd__a221o_1
X_8428_ _8231_/A _8231_/B _8230_/A _8333_/Y _8335_/A VGND VGND VPWR VPWR _8429_/B
+ sky130_fd_sc_hd__o311ai_4
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8359_ _8359_/A _8447_/B VGND VGND VPWR VPWR _8481_/B sky130_fd_sc_hd__or2_1
XFILLER_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5991_ _6041_/A _5991_/B VGND VGND VPWR VPWR _6037_/B sky130_fd_sc_hd__nor2_1
X_7730_ _7730_/A _7730_/B VGND VGND VPWR VPWR _7731_/B sky130_fd_sc_hd__nand2_1
X_4942_ _4943_/A _4943_/B VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7661_ _7661_/A _7661_/B _7660_/Y VGND VGND VPWR VPWR _7663_/A sky130_fd_sc_hd__nor3b_2
XFILLER_32_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6612_ _6710_/B _6612_/B VGND VGND VPWR VPWR _6614_/A sky130_fd_sc_hd__and2_1
X_4873_ _4873_/A VGND VGND VPWR VPWR _4873_/Y sky130_fd_sc_hd__clkinv_2
X_7592_ _7592_/A _7592_/B VGND VGND VPWR VPWR _7594_/B sky130_fd_sc_hd__xnor2_1
X_6543_ _6543_/A _6543_/B _6616_/A VGND VGND VPWR VPWR _6616_/B sky130_fd_sc_hd__nand3_2
X_6474_ _6480_/A _6480_/B _6560_/A VGND VGND VPWR VPWR _6475_/B sky130_fd_sc_hd__o21ai_1
X_8213_ _8850_/B VGND VGND VPWR VPWR _8898_/B sky130_fd_sc_hd__clkbuf_2
X_5425_ _5424_/X _5276_/X _5105_/A VGND VGND VPWR VPWR _5425_/Y sky130_fd_sc_hd__a21oi_1
X_9193_ _9213_/CLK _9193_/D VGND VGND VPWR VPWR _9193_/Q sky130_fd_sc_hd__dfxtp_1
X_8144_ _8144_/A _8144_/B VGND VGND VPWR VPWR _8145_/B sky130_fd_sc_hd__or2_1
X_5356_ _5200_/X _5355_/X _5575_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
X_8075_ _8137_/A _8351_/B VGND VGND VPWR VPWR _8076_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5287_ _5287_/A VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7026_ _7027_/B _7141_/A _7027_/A VGND VGND VPWR VPWR _7028_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8977_ _8974_/Y _9002_/B _8976_/X VGND VGND VPWR VPWR _8980_/A sky130_fd_sc_hd__o21a_1
XFILLER_82_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7928_ _8032_/A _8039_/A _7810_/D _7808_/X VGND VGND VPWR VPWR _7929_/B sky130_fd_sc_hd__a31o_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7859_ _7859_/A _7859_/B VGND VGND VPWR VPWR _7860_/B sky130_fd_sc_hd__and2_1
XFILLER_51_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5210_ _5210_/A VGND VGND VPWR VPWR _5653_/A sky130_fd_sc_hd__buf_2
XFILLER_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6190_ _7042_/D VGND VGND VPWR VPWR _6361_/D sky130_fd_sc_hd__buf_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5141_ _5141_/A VGND VGND VPWR VPWR _5151_/A sky130_fd_sc_hd__clkbuf_2
X_5072_ _5072_/A VGND VGND VPWR VPWR _5080_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8900_ _8900_/A _8900_/B VGND VGND VPWR VPWR _8945_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8831_ _8831_/A _8831_/B VGND VGND VPWR VPWR _8937_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8762_ _8761_/A _8761_/B _8760_/X VGND VGND VPWR VPWR _8825_/A sky130_fd_sc_hd__o21bai_1
X_7713_ _7830_/B _7713_/B VGND VGND VPWR VPWR _7716_/A sky130_fd_sc_hd__or2_1
X_5974_ _5974_/A _5974_/B VGND VGND VPWR VPWR _5976_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8693_ _8750_/A _8694_/C _8694_/A VGND VGND VPWR VPWR _8695_/A sky130_fd_sc_hd__a21oi_1
X_4925_ _4925_/A _4950_/B VGND VGND VPWR VPWR _4925_/Y sky130_fd_sc_hd__nor2_1
X_7644_ _7644_/A _7761_/A VGND VGND VPWR VPWR _7764_/A sky130_fd_sc_hd__nor2_1
X_4856_ _4856_/A _4856_/B VGND VGND VPWR VPWR _4856_/Y sky130_fd_sc_hd__nand2_1
X_7575_ _7576_/A _7576_/B VGND VGND VPWR VPWR _7577_/A sky130_fd_sc_hd__nor2_1
X_6526_ _7361_/C _7706_/A VGND VGND VPWR VPWR _6532_/A sky130_fd_sc_hd__nand2_1
X_4787_ _5621_/A _4787_/B VGND VGND VPWR VPWR _4787_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6457_ _6457_/A _6541_/B VGND VGND VPWR VPWR _6458_/C sky130_fd_sc_hd__nand2_2
X_9176_ _9216_/CLK input6/X VGND VGND VPWR VPWR _9176_/Q sky130_fd_sc_hd__dfxtp_1
X_6388_ _9205_/Q VGND VGND VPWR VPWR _7222_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5408_ _5368_/X _5581_/A _5406_/X _5407_/Y _5156_/X VGND VGND VPWR VPWR _5408_/X
+ sky130_fd_sc_hd__a221o_1
X_8127_ _8024_/A _8024_/B _8026_/Y _8019_/B _8126_/X VGND VGND VPWR VPWR _8231_/B
+ sky130_fd_sc_hd__a311oi_4
X_5339_ _5339_/A VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8058_ _8058_/A _8058_/B _8057_/X VGND VGND VPWR VPWR _8060_/A sky130_fd_sc_hd__or3b_1
XFILLER_75_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7009_ _7009_/A _7009_/B VGND VGND VPWR VPWR _7011_/A sky130_fd_sc_hd__xnor2_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X VGND VGND VPWR VPWR _9224_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5690_ _5160_/A _5689_/X _5734_/S VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__mux2_1
X_4710_ _9097_/Q VGND VGND VPWR VPWR _5728_/S sky130_fd_sc_hd__inv_2
X_4641_ _4641_/A VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__buf_2
X_7360_ _7360_/A VGND VGND VPWR VPWR _7756_/A sky130_fd_sc_hd__clkbuf_2
X_4572_ _4572_/A VGND VGND VPWR VPWR _4573_/A sky130_fd_sc_hd__clkbuf_2
X_6311_ _7019_/C VGND VGND VPWR VPWR _7129_/B sky130_fd_sc_hd__clkbuf_2
X_7291_ _6974_/B _9211_/Q _9212_/Q _6974_/A VGND VGND VPWR VPWR _7295_/D sky130_fd_sc_hd__a22o_1
X_9030_ _9029_/A _9029_/B _9029_/C VGND VGND VPWR VPWR _9031_/B sky130_fd_sc_hd__a21oi_1
X_6242_ _6342_/A _6242_/B VGND VGND VPWR VPWR _6335_/B sky130_fd_sc_hd__or2_1
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6173_ _6974_/A VGND VGND VPWR VPWR _6251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5124_ _5124_/A VGND VGND VPWR VPWR _5124_/X sky130_fd_sc_hd__buf_2
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5055_ _5051_/Y _5054_/X _5154_/A VGND VGND VPWR VPWR _5055_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8814_ _8814_/A _8814_/B VGND VGND VPWR VPWR _8815_/B sky130_fd_sc_hd__or2_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8745_ _8745_/A _8688_/C VGND VGND VPWR VPWR _8746_/C sky130_fd_sc_hd__or2b_1
X_5957_ _9052_/B _5957_/B VGND VGND VPWR VPWR _5958_/A sky130_fd_sc_hd__and2_1
XFILLER_40_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8676_ _8909_/A _8844_/A _8844_/C _8867_/A VGND VGND VPWR VPWR _8678_/A sky130_fd_sc_hd__a22oi_2
X_4908_ _4939_/B VGND VGND VPWR VPWR _4937_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7627_ _7627_/A _8091_/C VGND VGND VPWR VPWR _7754_/A sky130_fd_sc_hd__nand2_1
X_5888_ _6022_/A _7253_/A VGND VGND VPWR VPWR _5987_/A sky130_fd_sc_hd__nand2_2
X_4839_ _4839_/A VGND VGND VPWR VPWR _5215_/A sky130_fd_sc_hd__clkbuf_2
X_7558_ _7425_/A _7425_/B _7429_/B VGND VGND VPWR VPWR _7558_/Y sky130_fd_sc_hd__a21oi_1
X_7489_ _7628_/A _7756_/A VGND VGND VPWR VPWR _7490_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _6508_/A _6508_/B _6508_/C VGND VGND VPWR VPWR _6637_/A sky130_fd_sc_hd__a21o_1
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9159_ _9214_/CLK _9159_/D VGND VGND VPWR VPWR _9159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A VGND VGND VPWR VPWR clkbuf_4_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_6 _9068_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6860_ _6251_/A _7706_/C _7583_/D _6825_/A VGND VGND VPWR VPWR _6861_/B sky130_fd_sc_hd__a22oi_1
X_6791_ _6791_/A _6791_/B VGND VGND VPWR VPWR _6793_/A sky130_fd_sc_hd__xnor2_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5811_ _5940_/A _5809_/X _5810_/X VGND VGND VPWR VPWR _5812_/B sky130_fd_sc_hd__a21bo_1
X_8530_ _8530_/A _8538_/A _8792_/B _8733_/D VGND VGND VPWR VPWR _8530_/X sky130_fd_sc_hd__and4_1
X_5742_ _4889_/X _5741_/X _5742_/S VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__mux2_1
X_8461_ _8597_/A VGND VGND VPWR VPWR _8756_/A sky130_fd_sc_hd__buf_2
X_5673_ _5754_/A _5672_/X _5673_/S VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8392_ _8392_/A _8392_/B VGND VGND VPWR VPWR _8392_/Y sky130_fd_sc_hd__xnor2_1
X_4624_ _5697_/S VGND VGND VPWR VPWR _5282_/S sky130_fd_sc_hd__clkbuf_2
X_7412_ _9215_/Q VGND VGND VPWR VPWR _7804_/B sky130_fd_sc_hd__clkbuf_2
X_7343_ _7340_/X _7341_/Y _7342_/X _7234_/B VGND VGND VPWR VPWR _7380_/A sky130_fd_sc_hd__o211a_1
X_4555_ _5000_/A VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9013_ _9013_/A _9013_/B VGND VGND VPWR VPWR _9035_/A sky130_fd_sc_hd__or2_1
X_7274_ _7274_/A _7274_/B _7274_/C VGND VGND VPWR VPWR _7277_/C sky130_fd_sc_hd__and3_1
X_6225_ _7509_/A _7457_/A _6329_/A _6228_/D VGND VGND VPWR VPWR _6231_/A sky130_fd_sc_hd__a22o_1
XFILLER_97_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6156_ _6922_/B _6313_/B _7457_/A _6313_/A VGND VGND VPWR VPWR _6157_/B sky130_fd_sc_hd__a22oi_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _4891_/A _5106_/X _5095_/X VGND VGND VPWR VPWR _5107_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6087_ _6087_/A _6087_/B _6087_/C VGND VGND VPWR VPWR _6090_/B sky130_fd_sc_hd__nand3_1
XFILLER_26_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5038_ _5074_/B VGND VGND VPWR VPWR _5080_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8728_ _8727_/B _8728_/B VGND VGND VPWR VPWR _8729_/B sky130_fd_sc_hd__and2b_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6989_ _6988_/A _6988_/B _6988_/C VGND VGND VPWR VPWR _7174_/A sky130_fd_sc_hd__a21oi_1
XFILLER_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8659_ _8716_/A _9025_/A _9029_/B _8438_/B VGND VGND VPWR VPWR _8691_/A sky130_fd_sc_hd__a22oi_1
XFILLER_21_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput76 _9130_/Q VGND VGND VPWR VPWR F[1] sky130_fd_sc_hd__buf_2
Xoutput65 _9129_/Q VGND VGND VPWR VPWR F[0] sky130_fd_sc_hd__buf_2
Xoutput87 _9131_/Q VGND VGND VPWR VPWR F[2] sky130_fd_sc_hd__buf_2
XFILLER_76_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6010_ _6010_/A _6010_/B _6010_/C VGND VGND VPWR VPWR _6018_/C sky130_fd_sc_hd__nand3_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7961_ _8190_/A VGND VGND VPWR VPWR _8379_/A sky130_fd_sc_hd__buf_2
XFILLER_67_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7892_ _7891_/A _7891_/B _7891_/C VGND VGND VPWR VPWR _7893_/B sky130_fd_sc_hd__a21o_1
X_6912_ _6913_/B _7029_/A _6913_/A VGND VGND VPWR VPWR _6912_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ _6843_/A _6843_/B _6843_/C VGND VGND VPWR VPWR _6844_/B sky130_fd_sc_hd__and3_1
X_6774_ _6774_/A _6774_/B VGND VGND VPWR VPWR _6795_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8513_ _8513_/A _8513_/B VGND VGND VPWR VPWR _8513_/Y sky130_fd_sc_hd__nor2_1
X_5725_ _9091_/Q _4568_/A _5724_/X _4857_/A VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__o211a_1
X_8444_ _8444_/A _8444_/B VGND VGND VPWR VPWR _8525_/B sky130_fd_sc_hd__nand2_1
X_5656_ _5656_/A _5656_/B VGND VGND VPWR VPWR _5656_/Y sky130_fd_sc_hd__nand2_1
X_4607_ _4607_/A VGND VGND VPWR VPWR _4637_/A sky130_fd_sc_hd__clkbuf_2
X_8375_ _8492_/B _8375_/B VGND VGND VPWR VPWR _8377_/A sky130_fd_sc_hd__xnor2_1
X_5587_ _5251_/A _9086_/Q _5585_/X _5586_/X _4786_/S VGND VGND VPWR VPWR _5587_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7326_ _7042_/C _7327_/C _7148_/D _7153_/C VGND VGND VPWR VPWR _7328_/A sky130_fd_sc_hd__a22oi_1
X_4538_ _4538_/A VGND VGND VPWR VPWR _5765_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7257_ _7257_/A _7640_/A VGND VGND VPWR VPWR _7261_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6208_ _6118_/A _6118_/B _6118_/C VGND VGND VPWR VPWR _6210_/C sky130_fd_sc_hd__a21bo_1
XFILLER_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7188_ _6968_/A _7571_/A _7186_/Y _7187_/X VGND VGND VPWR VPWR _7190_/A sky130_fd_sc_hd__o2bb2a_1
X_6139_ _6139_/A VGND VGND VPWR VPWR _6325_/A sky130_fd_sc_hd__clkbuf_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5510_ _5510_/A VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__buf_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6490_ _6859_/B VGND VGND VPWR VPWR _7187_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ _5247_/X _5273_/X _5378_/X VGND VGND VPWR VPWR _5441_/Y sky130_fd_sc_hd__a21oi_1
X_8160_ _8092_/A _8094_/B _8092_/B VGND VGND VPWR VPWR _8161_/B sky130_fd_sc_hd__o21ba_1
X_5372_ _5558_/A _5482_/A _4676_/C _5430_/A _4572_/A VGND VGND VPWR VPWR _5372_/X
+ sky130_fd_sc_hd__o221a_1
X_8091_ _8091_/A _8091_/B _8091_/C _8091_/D VGND VGND VPWR VPWR _8092_/B sky130_fd_sc_hd__and4_1
X_7111_ _9197_/Q _9182_/Q VGND VGND VPWR VPWR _7767_/C sky130_fd_sc_hd__and2_2
XFILLER_99_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7042_ _7327_/A _7042_/B _7042_/C _7042_/D VGND VGND VPWR VPWR _7043_/B sky130_fd_sc_hd__and4_1
XFILLER_101_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8993_ _9013_/A _8994_/C _8954_/A _8954_/B VGND VGND VPWR VPWR _8993_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7944_ _7944_/A _7944_/B _7944_/C VGND VGND VPWR VPWR _7945_/B sky130_fd_sc_hd__nor3_1
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7875_ _7876_/A _7876_/B VGND VGND VPWR VPWR _7877_/A sky130_fd_sc_hd__or2_1
XFILLER_82_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6826_ _6831_/B _6822_/Y _6825_/X VGND VGND VPWR VPWR _6829_/A sky130_fd_sc_hd__a21oi_4
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6757_ _6757_/A _6757_/B VGND VGND VPWR VPWR _6766_/A sky130_fd_sc_hd__xnor2_2
X_5708_ _5618_/X _5136_/X _5367_/A VGND VGND VPWR VPWR _5708_/Y sky130_fd_sc_hd__a21oi_1
X_6688_ _6689_/B _6810_/A _6689_/A VGND VGND VPWR VPWR _6690_/A sky130_fd_sc_hd__a21o_1
X_8427_ _8510_/B _8427_/B VGND VGND VPWR VPWR _8430_/A sky130_fd_sc_hd__nor2_1
X_5639_ _5394_/A _5249_/X _4667_/A VGND VGND VPWR VPWR _5639_/Y sky130_fd_sc_hd__a21oi_1
X_8358_ _8358_/A _8358_/B VGND VGND VPWR VPWR _8447_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7309_ _7309_/A _7309_/B VGND VGND VPWR VPWR _7310_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8289_ _8607_/B VGND VGND VPWR VPWR _8664_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5990_ _5989_/B _5990_/B VGND VGND VPWR VPWR _5991_/B sky130_fd_sc_hd__and2b_1
XFILLER_64_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ _5146_/A _4936_/Y _4937_/X _4940_/X VGND VGND VPWR VPWR _4941_/X sky130_fd_sc_hd__a31o_1
X_7660_ _7660_/A _7660_/B VGND VGND VPWR VPWR _7660_/Y sky130_fd_sc_hd__xnor2_1
X_4872_ _4850_/B _4870_/X _4872_/S VGND VGND VPWR VPWR _4872_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6611_ _6611_/A _6611_/B _6611_/C VGND VGND VPWR VPWR _6612_/B sky130_fd_sc_hd__or3_1
X_7591_ _7440_/A _7440_/B _7590_/X VGND VGND VPWR VPWR _7592_/B sky130_fd_sc_hd__a21oi_1
X_6542_ _6541_/A _6541_/B _6541_/C VGND VGND VPWR VPWR _6616_/A sky130_fd_sc_hd__a21o_1
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6473_ _6473_/A _6379_/B VGND VGND VPWR VPWR _6560_/A sky130_fd_sc_hd__or2b_1
X_8212_ _8211_/A _8211_/B _8211_/C VGND VGND VPWR VPWR _8223_/C sky130_fd_sc_hd__a21oi_2
X_9192_ _9216_/CLK _9192_/D VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
X_5424_ _5424_/A VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__buf_2
X_8143_ _8144_/A _8144_/B VGND VGND VPWR VPWR _8254_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5355_ _5117_/A _5354_/X _5527_/S VGND VGND VPWR VPWR _5355_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8074_ _8664_/D VGND VGND VPWR VPWR _8351_/B sky130_fd_sc_hd__clkbuf_2
X_5286_ _5286_/A VGND VGND VPWR VPWR _5287_/A sky130_fd_sc_hd__buf_2
X_7025_ _7145_/A _7025_/B VGND VGND VPWR VPWR _7027_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8976_ _8975_/A _8891_/B _8978_/B _8974_/A VGND VGND VPWR VPWR _8976_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7927_ _7927_/A _7927_/B VGND VGND VPWR VPWR _7929_/A sky130_fd_sc_hd__xnor2_1
X_7858_ _7859_/A _7859_/B VGND VGND VPWR VPWR _7860_/A sky130_fd_sc_hd__nor2_1
X_6809_ _6809_/A _6809_/B VGND VGND VPWR VPWR _6810_/C sky130_fd_sc_hd__nand2_2
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7789_ _7788_/A _7788_/B _7788_/C VGND VGND VPWR VPWR _7790_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5140_ _5140_/A VGND VGND VPWR VPWR _5141_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5071_ _5071_/A VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8830_ _8830_/A _8818_/B VGND VGND VPWR VPWR _8872_/B sky130_fd_sc_hd__or2b_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8761_ _8761_/A _8761_/B _8760_/X VGND VGND VPWR VPWR _8763_/A sky130_fd_sc_hd__or3b_1
X_5973_ _6859_/B _7254_/C VGND VGND VPWR VPWR _5974_/B sky130_fd_sc_hd__nand2_1
X_7712_ _7712_/A _7712_/B _7712_/C VGND VGND VPWR VPWR _7713_/B sky130_fd_sc_hd__nor3_1
X_4924_ _4924_/A _4950_/A VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__or2_1
X_8692_ _8691_/A _8726_/A _8691_/C _8753_/B VGND VGND VPWR VPWR _8694_/C sky130_fd_sc_hd__o22ai_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7643_ _7643_/A _7643_/B VGND VGND VPWR VPWR _7761_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4855_ _5144_/A _4830_/X _4850_/Y _4854_/X VGND VGND VPWR VPWR _4855_/X sky130_fd_sc_hd__o2bb2a_1
X_7574_ _7689_/A _9214_/Q VGND VGND VPWR VPWR _7576_/B sky130_fd_sc_hd__and2_1
X_4786_ _4760_/X _4785_/X _4786_/S VGND VGND VPWR VPWR _4786_/X sky130_fd_sc_hd__mux2_1
X_6525_ _6525_/A _6454_/A VGND VGND VPWR VPWR _6541_/A sky130_fd_sc_hd__or2b_1
X_6456_ _6456_/A _6456_/B VGND VGND VPWR VPWR _6541_/B sky130_fd_sc_hd__nand2_1
X_9175_ _9210_/CLK input5/X VGND VGND VPWR VPWR _9175_/Q sky130_fd_sc_hd__dfxtp_2
X_5407_ _5142_/X _5485_/A _5154_/X VGND VGND VPWR VPWR _5407_/Y sky130_fd_sc_hd__a21oi_1
X_6387_ _6345_/A _6387_/B VGND VGND VPWR VPWR _6411_/B sky130_fd_sc_hd__and2b_1
X_8126_ _8231_/A _8126_/B VGND VGND VPWR VPWR _8126_/X sky130_fd_sc_hd__or2_1
X_5338_ _5315_/X _5202_/X _5204_/X _5336_/X _5337_/X VGND VGND VPWR VPWR _9133_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8057_ _8197_/B _8057_/B VGND VGND VPWR VPWR _8057_/X sky130_fd_sc_hd__or2_1
X_7008_ _7008_/A _7008_/B VGND VGND VPWR VPWR _7009_/B sky130_fd_sc_hd__nor2_1
X_5269_ _5129_/X _5212_/X _5265_/X _5268_/Y _5175_/X VGND VGND VPWR VPWR _5269_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8959_ _8959_/A _8959_/B VGND VGND VPWR VPWR _8959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4640_ _5071_/A VGND VGND VPWR VPWR _4641_/A sky130_fd_sc_hd__clkbuf_2
X_6310_ _9174_/Q VGND VGND VPWR VPWR _7019_/C sky130_fd_sc_hd__clkbuf_2
X_4571_ _4571_/A VGND VGND VPWR VPWR _4572_/A sky130_fd_sc_hd__clkbuf_2
X_7290_ _7290_/A _7552_/B VGND VGND VPWR VPWR _9088_/D sky130_fd_sc_hd__xor2_1
XFILLER_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6241_ _6778_/B _6925_/A _7455_/A _6886_/A VGND VGND VPWR VPWR _6242_/B sky130_fd_sc_hd__a22oi_4
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6172_ _6172_/A VGND VGND VPWR VPWR _6907_/A sky130_fd_sc_hd__buf_2
XFILLER_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _9084_/Q VGND VGND VPWR VPWR _5124_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5054_ _5053_/A _5053_/Y _5054_/S VGND VGND VPWR VPWR _5054_/X sky130_fd_sc_hd__mux2_1
X_8813_ _8814_/A _8814_/B VGND VGND VPWR VPWR _8813_/X sky130_fd_sc_hd__and2_1
XFILLER_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8744_ _8744_/A _8744_/B VGND VGND VPWR VPWR _8806_/B sky130_fd_sc_hd__or2_1
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5956_ _9052_/A _5954_/B _9055_/A VGND VGND VPWR VPWR _5957_/B sky130_fd_sc_hd__a21o_1
X_5887_ _9193_/Q VGND VGND VPWR VPWR _7253_/A sky130_fd_sc_hd__buf_2
X_8675_ _8675_/A VGND VGND VPWR VPWR _8867_/A sky130_fd_sc_hd__clkbuf_2
X_4907_ _4913_/A _4913_/B VGND VGND VPWR VPWR _4939_/B sky130_fd_sc_hd__xor2_2
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7626_ _8137_/A _8595_/A _7492_/B _7490_/Y VGND VGND VPWR VPWR _7637_/A sky130_fd_sc_hd__a31o_1
X_4838_ _4927_/A _4963_/A VGND VGND VPWR VPWR _4838_/Y sky130_fd_sc_hd__nor2_4
X_4769_ _4769_/A _4769_/B VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__nand2_1
X_7557_ _7531_/A _8756_/B _7536_/B _7535_/B VGND VGND VPWR VPWR _7672_/A sky130_fd_sc_hd__a31o_1
X_7488_ _7627_/A _7756_/A VGND VGND VPWR VPWR _7629_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6508_ _6508_/A _6508_/B _6508_/C VGND VGND VPWR VPWR _6508_/X sky130_fd_sc_hd__and3_1
X_6439_ _6313_/B _7583_/B _7728_/C _6313_/A VGND VGND VPWR VPWR _6444_/A sky130_fd_sc_hd__a22oi_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9158_ _9199_/CLK _9158_/D VGND VGND VPWR VPWR _9158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8109_ _8135_/A _8135_/B VGND VGND VPWR VPWR _8111_/C sky130_fd_sc_hd__xnor2_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_9089_ _9090_/CLK _9089_/D VGND VGND VPWR VPWR _9089_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_7 _9075_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6790_ _6790_/A _6790_/B VGND VGND VPWR VPWR _6791_/B sky130_fd_sc_hd__nor2_1
X_5810_ _7367_/B _6025_/A _9163_/Q _7367_/A VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5741_ _4541_/A _5740_/X _5741_/S VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__mux2_1
X_8460_ _8460_/A _8460_/B VGND VGND VPWR VPWR _8480_/A sky130_fd_sc_hd__xor2_1
X_5672_ _5557_/A _5671_/X _5695_/S VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__mux2_1
X_7411_ _7411_/A VGND VGND VPWR VPWR _7544_/B sky130_fd_sc_hd__inv_2
X_8391_ _8391_/A _8474_/B VGND VGND VPWR VPWR _8392_/B sky130_fd_sc_hd__xnor2_1
X_4623_ _5741_/S VGND VGND VPWR VPWR _5697_/S sky130_fd_sc_hd__clkbuf_2
X_7342_ _7342_/A _7342_/B _7342_/C VGND VGND VPWR VPWR _7342_/X sky130_fd_sc_hd__or3_1
X_4554_ _9100_/Q VGND VGND VPWR VPWR _5000_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7273_ _7383_/B _7273_/B VGND VGND VPWR VPWR _7274_/C sky130_fd_sc_hd__nand2_2
X_9012_ _9013_/A _9013_/B VGND VGND VPWR VPWR _9014_/A sky130_fd_sc_hd__nand2_1
X_6224_ _6325_/A _7148_/B _6143_/B _6325_/B VGND VGND VPWR VPWR _6228_/D sky130_fd_sc_hd__a22o_1
X_6155_ _7042_/C VGND VGND VPWR VPWR _7457_/A sky130_fd_sc_hd__clkbuf_4
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6086_ _6087_/B _6087_/C _6087_/A VGND VGND VPWR VPWR _6090_/A sky130_fd_sc_hd__a21o_1
X_5106_ _5089_/X _5105_/Y _5090_/X VGND VGND VPWR VPWR _5106_/X sky130_fd_sc_hd__o21a_1
X_5037_ _5067_/B VGND VGND VPWR VPWR _5074_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8727_ _8728_/B _8727_/B VGND VGND VPWR VPWR _8729_/A sky130_fd_sc_hd__and2b_1
X_6988_ _6988_/A _6988_/B _6988_/C VGND VGND VPWR VPWR _6988_/X sky130_fd_sc_hd__and3_1
XFILLER_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5939_ _5987_/A _5939_/B VGND VGND VPWR VPWR _5948_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8658_ _8978_/B VGND VGND VPWR VPWR _9029_/B sky130_fd_sc_hd__clkbuf_2
X_8589_ _8586_/Y _8668_/A _8716_/A _8844_/D VGND VGND VPWR VPWR _8668_/B sky130_fd_sc_hd__and4bb_1
X_7609_ _8243_/A _7847_/D _7959_/D _7852_/A VGND VGND VPWR VPWR _7611_/A sky130_fd_sc_hd__a22oi_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X VGND VGND VPWR VPWR _9220_/CLK sky130_fd_sc_hd__clkbuf_2
Xoutput66 _9139_/Q VGND VGND VPWR VPWR F[10] sky130_fd_sc_hd__buf_2
Xoutput77 _9149_/Q VGND VGND VPWR VPWR F[20] sky130_fd_sc_hd__buf_2
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput88 _9159_/Q VGND VGND VPWR VPWR F[30] sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7960_ _7960_/A _7960_/B VGND VGND VPWR VPWR _7963_/A sky130_fd_sc_hd__nor2_1
X_7891_ _7891_/A _7891_/B _7891_/C VGND VGND VPWR VPWR _7893_/A sky130_fd_sc_hd__nand3_1
X_6911_ _7034_/A _6911_/B VGND VGND VPWR VPWR _6913_/A sky130_fd_sc_hd__xnor2_2
XFILLER_35_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6842_ _6843_/B _6843_/C _6843_/A VGND VGND VPWR VPWR _6844_/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6773_ _6773_/A _6673_/A VGND VGND VPWR VPWR _6795_/A sky130_fd_sc_hd__or2b_1
X_8512_ _8512_/A _8512_/B VGND VGND VPWR VPWR _9099_/D sky130_fd_sc_hd__xor2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5724_ _9089_/Q _4778_/A _5723_/X _9094_/Q VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a211o_1
X_8443_ _8444_/A _8444_/B VGND VGND VPWR VPWR _8445_/A sky130_fd_sc_hd__or2_1
X_5655_ _5734_/S VGND VGND VPWR VPWR _5712_/S sky130_fd_sc_hd__clkbuf_2
X_8374_ _8278_/A _8282_/B _8278_/B VGND VGND VPWR VPWR _8375_/B sky130_fd_sc_hd__o21ba_1
X_4606_ _5132_/A VGND VGND VPWR VPWR _4607_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7325_ _7325_/A _9207_/Q VGND VGND VPWR VPWR _7329_/A sky130_fd_sc_hd__nand2_1
X_5586_ _4856_/A _5208_/A _5141_/A VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4537_ _4737_/A VGND VGND VPWR VPWR _4538_/A sky130_fd_sc_hd__clkbuf_2
X_7256_ _7352_/B _7256_/B VGND VGND VPWR VPWR _7357_/A sky130_fd_sc_hd__nor2_1
X_6207_ _6207_/A _6207_/B _6207_/C VGND VGND VPWR VPWR _6210_/B sky130_fd_sc_hd__nand3_1
X_7187_ _7187_/A _7187_/B _7694_/C _7694_/D VGND VGND VPWR VPWR _7187_/X sky130_fd_sc_hd__and4_1
X_6138_ _7770_/A _6223_/B _6607_/A _7040_/A VGND VGND VPWR VPWR _6145_/B sky130_fd_sc_hd__nand4_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6069_ _6007_/A _6007_/C _6007_/B VGND VGND VPWR VPWR _6071_/C sky130_fd_sc_hd__a21bo_1
XFILLER_73_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5440_ _5160_/X _5653_/A _5438_/X _5439_/Y _5410_/X VGND VGND VPWR VPWR _5440_/X
+ sky130_fd_sc_hd__a221o_1
X_5371_ _5371_/A VGND VGND VPWR VPWR _5558_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8090_ _8156_/B _7966_/D _8091_/D _8154_/A VGND VGND VPWR VPWR _8092_/A sky130_fd_sc_hd__a22oi_1
X_7110_ _7110_/A _7110_/B VGND VGND VPWR VPWR _7126_/B sky130_fd_sc_hd__nand2_1
X_7041_ _6759_/C _7822_/A _6572_/D _6143_/B VGND VGND VPWR VPWR _7043_/A sky130_fd_sc_hd__a22oi_1
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8992_ _8992_/A _8992_/B VGND VGND VPWR VPWR _8994_/C sky130_fd_sc_hd__nand2_1
XFILLER_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7943_ _7944_/A _7944_/B _7944_/C VGND VGND VPWR VPWR _8058_/B sky130_fd_sc_hd__o21a_1
X_7874_ _7874_/A _7874_/B VGND VGND VPWR VPWR _7876_/B sky130_fd_sc_hd__xnor2_1
X_6825_ _6825_/A _6825_/B _6825_/C _7822_/D VGND VGND VPWR VPWR _6825_/X sky130_fd_sc_hd__and4_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6756_ _6756_/A _6756_/B VGND VGND VPWR VPWR _6757_/B sky130_fd_sc_hd__nor2_1
X_5707_ _4650_/A _5258_/X _5705_/X _5706_/Y _4599_/A VGND VGND VPWR VPWR _5707_/X
+ sky130_fd_sc_hd__a221o_1
X_6687_ _6752_/A _6687_/B VGND VGND VPWR VPWR _6689_/A sky130_fd_sc_hd__xnor2_1
XFILLER_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8426_ _8423_/Y _8424_/X _8328_/B _8336_/X VGND VGND VPWR VPWR _8427_/B sky130_fd_sc_hd__o211a_1
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5638_ _4634_/A _5116_/A _5636_/X _5637_/Y _5249_/X VGND VGND VPWR VPWR _5638_/X
+ sky130_fd_sc_hd__a221o_1
X_8357_ _8358_/A _8358_/B VGND VGND VPWR VPWR _8359_/A sky130_fd_sc_hd__and2_1
X_5569_ _5287_/A _4723_/X _4672_/A VGND VGND VPWR VPWR _5569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7308_ _7308_/A _7308_/B VGND VGND VPWR VPWR _7310_/A sky130_fd_sc_hd__nor2_1
X_8288_ _8721_/A VGND VGND VPWR VPWR _8664_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7239_ _7237_/X _7160_/B _7235_/Y _7319_/A VGND VGND VPWR VPWR _7319_/B sky130_fd_sc_hd__o211ai_4
XFILLER_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4940_ _4940_/A _4940_/B _4940_/C VGND VGND VPWR VPWR _4940_/X sky130_fd_sc_hd__and3_1
XFILLER_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4871_ _5730_/S VGND VGND VPWR VPWR _4872_/S sky130_fd_sc_hd__buf_2
X_7590_ _7439_/A _7590_/B VGND VGND VPWR VPWR _7590_/X sky130_fd_sc_hd__and2b_1
XFILLER_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6610_ _6611_/A _6611_/B _6611_/C VGND VGND VPWR VPWR _6710_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6541_ _6541_/A _6541_/B _6541_/C VGND VGND VPWR VPWR _6543_/B sky130_fd_sc_hd__nand3_1
X_6472_ _6481_/A _6481_/B VGND VGND VPWR VPWR _6560_/B sky130_fd_sc_hd__xnor2_2
X_8211_ _8211_/A _8211_/B _8211_/C VGND VGND VPWR VPWR _8223_/B sky130_fd_sc_hd__and3_1
X_5423_ _9091_/Q VGND VGND VPWR VPWR _5424_/A sky130_fd_sc_hd__inv_2
X_9191_ _9216_/CLK _9191_/D VGND VGND VPWR VPWR _9191_/Q sky130_fd_sc_hd__dfxtp_4
X_8142_ _7747_/X _8844_/D _8076_/A _8072_/B VGND VGND VPWR VPWR _8144_/B sky130_fd_sc_hd__a31o_1
X_5354_ _5120_/A _5353_/X _5354_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8073_ _8721_/B VGND VGND VPWR VPWR _8664_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5285_ _5245_/X _5202_/X _5204_/X _5283_/X _5284_/X VGND VGND VPWR VPWR _9131_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7024_ _7024_/A _7161_/A VGND VGND VPWR VPWR _7025_/B sky130_fd_sc_hd__and2_1
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8975_ _8975_/A _8978_/B VGND VGND VPWR VPWR _9002_/B sky130_fd_sc_hd__nand2_1
X_7926_ _8220_/A _8039_/A VGND VGND VPWR VPWR _7927_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7857_ _7978_/B _7857_/B VGND VGND VPWR VPWR _7859_/B sky130_fd_sc_hd__xnor2_1
X_6808_ _6808_/A _6808_/B _6808_/C VGND VGND VPWR VPWR _6809_/B sky130_fd_sc_hd__nand3_2
XFILLER_51_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7788_ _7788_/A _7788_/B _7788_/C VGND VGND VPWR VPWR _7790_/A sky130_fd_sc_hd__and3_1
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _6740_/B _6740_/C _6740_/A VGND VGND VPWR VPWR _6845_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8409_ _8981_/B VGND VGND VPWR VPWR _9029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5070_ _5063_/Y _5066_/X _5069_/X _4875_/S _5733_/S VGND VGND VPWR VPWR _5070_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_49_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8760_ _8760_/A _8819_/B VGND VGND VPWR VPWR _8760_/X sky130_fd_sc_hd__or2_1
X_5972_ _9198_/Q VGND VGND VPWR VPWR _7254_/C sky130_fd_sc_hd__buf_2
X_7711_ _7712_/A _7712_/B _7712_/C VGND VGND VPWR VPWR _7830_/B sky130_fd_sc_hd__o21a_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4923_ _4923_/A VGND VGND VPWR VPWR _5382_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8691_ _8691_/A _8726_/A _8691_/C _8753_/B VGND VGND VPWR VPWR _8750_/A sky130_fd_sc_hd__or4_4
X_7642_ _7880_/A _8721_/B VGND VGND VPWR VPWR _7643_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _5286_/A _4873_/A _5144_/A VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__a21o_1
X_7573_ _7573_/A _7573_/B VGND VGND VPWR VPWR _7576_/A sky130_fd_sc_hd__xor2_1
X_4785_ _5140_/A _4764_/X _4782_/X _4784_/Y VGND VGND VPWR VPWR _4785_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6524_ _6566_/A _6524_/B VGND VGND VPWR VPWR _6543_/A sky130_fd_sc_hd__xnor2_1
X_6455_ _6456_/A _6456_/B VGND VGND VPWR VPWR _6457_/A sky130_fd_sc_hd__or2_1
X_9174_ _9210_/CLK input4/X VGND VGND VPWR VPWR _9174_/Q sky130_fd_sc_hd__dfxtp_2
X_5406_ _5149_/X _5532_/A _5404_/Y _5405_/X _5151_/X VGND VGND VPWR VPWR _5406_/X
+ sky130_fd_sc_hd__a221o_1
X_6386_ _6370_/A _6370_/B _6369_/B VGND VGND VPWR VPWR _6470_/A sky130_fd_sc_hd__a21o_1
XFILLER_87_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8125_ _8125_/A _8125_/B VGND VGND VPWR VPWR _8126_/B sky130_fd_sc_hd__and2_1
X_5337_ _9071_/Q _5337_/B VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__or2_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8056_ _8056_/A _8056_/B _8056_/C VGND VGND VPWR VPWR _8057_/B sky130_fd_sc_hd__nor3_1
X_5268_ _5266_/X _5604_/A _5173_/X VGND VGND VPWR VPWR _5268_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7007_ _6325_/A _7254_/D _7360_/A _6325_/B VGND VGND VPWR VPWR _7008_/B sky130_fd_sc_hd__a22oi_2
X_5199_ _5199_/A VGND VGND VPWR VPWR _9129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8958_ _8958_/A _8958_/B VGND VGND VPWR VPWR _8961_/A sky130_fd_sc_hd__or2_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7909_ _7796_/A _7796_/B _7792_/Y _7794_/B VGND VGND VPWR VPWR _7910_/B sky130_fd_sc_hd__o31a_1
X_8889_ _8889_/A _8889_/B VGND VGND VPWR VPWR _8890_/B sky130_fd_sc_hd__or2_1
XFILLER_70_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _4570_/A VGND VGND VPWR VPWR _4571_/A sky130_fd_sc_hd__clkbuf_2
X_6240_ _6240_/A VGND VGND VPWR VPWR _6886_/A sky130_fd_sc_hd__buf_2
X_6171_ _6859_/A _7083_/A _6257_/C _6907_/B VGND VGND VPWR VPWR _6175_/A sky130_fd_sc_hd__and4_1
X_5122_ _5122_/A VGND VGND VPWR VPWR _5122_/X sky130_fd_sc_hd__buf_2
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5053_ _5053_/A _5053_/B VGND VGND VPWR VPWR _5053_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8812_ _8812_/A _8812_/B VGND VGND VPWR VPWR _8814_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8743_ _8744_/A _8744_/B VGND VGND VPWR VPWR _8746_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5955_ _6126_/A VGND VGND VPWR VPWR _9052_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8674_ _8674_/A VGND VGND VPWR VPWR _8909_/A sky130_fd_sc_hd__buf_2
XFILLER_80_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ _4816_/A _4817_/S _4816_/B VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__a21oi_4
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5886_ _5886_/A _5886_/B VGND VGND VPWR VPWR _9059_/A sky130_fd_sc_hd__xor2_1
X_7625_ _8466_/A VGND VGND VPWR VPWR _8595_/A sky130_fd_sc_hd__buf_2
XFILLER_21_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4837_ _4837_/A _5074_/A VGND VGND VPWR VPWR _4963_/A sky130_fd_sc_hd__and2_2
XFILLER_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7556_ _8909_/B VGND VGND VPWR VPWR _8756_/B sky130_fd_sc_hd__clkbuf_4
X_4768_ _4852_/A _4866_/A VGND VGND VPWR VPWR _4769_/B sky130_fd_sc_hd__nor2_2
X_7487_ _8069_/A _7852_/C VGND VGND VPWR VPWR _7487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6507_ _6507_/A _6507_/B VGND VGND VPWR VPWR _6508_/C sky130_fd_sc_hd__xnor2_2
X_4699_ _5103_/A VGND VGND VPWR VPWR _5187_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6438_ _7241_/B VGND VGND VPWR VPWR _7728_/C sky130_fd_sc_hd__clkbuf_4
X_9157_ _9223_/CLK _9157_/D VGND VGND VPWR VPWR _9157_/Q sky130_fd_sc_hd__dfxtp_1
X_8108_ _7981_/A _8064_/B _8003_/B _8002_/B VGND VGND VPWR VPWR _8135_/B sky130_fd_sc_hd__a31o_1
X_6369_ _6369_/A _6369_/B VGND VGND VPWR VPWR _6370_/B sky130_fd_sc_hd__nor2_1
XFILLER_102_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_9088_ _9090_/CLK _9088_/D VGND VGND VPWR VPWR _9088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8039_ _8039_/A VGND VGND VPWR VPWR _8597_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_75_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_8 _9140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5740_ _5678_/A _5739_/X _5740_/S VGND VGND VPWR VPWR _5740_/X sky130_fd_sc_hd__mux2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7410_/A _7548_/B VGND VGND VPWR VPWR _9089_/D sky130_fd_sc_hd__nor2_1
X_5671_ _5534_/A _5670_/X _5671_/S VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__mux2_1
X_8390_ _8390_/A _8390_/B VGND VGND VPWR VPWR _8474_/B sky130_fd_sc_hd__xnor2_1
X_4622_ _9110_/Q VGND VGND VPWR VPWR _5741_/S sky130_fd_sc_hd__inv_2
X_7341_ _7340_/A _7340_/B _7340_/C VGND VGND VPWR VPWR _7341_/Y sky130_fd_sc_hd__a21oi_1
X_4553_ _5733_/S VGND VGND VPWR VPWR _4876_/A sky130_fd_sc_hd__buf_2
X_7272_ _7271_/A _7319_/B _7271_/C _7383_/A VGND VGND VPWR VPWR _7273_/B sky130_fd_sc_hd__a22o_1
X_9011_ _9032_/A _9011_/B VGND VGND VPWR VPWR _9013_/B sky130_fd_sc_hd__or2_1
X_6223_ _6223_/A _6223_/B _7040_/A _7453_/A VGND VGND VPWR VPWR _6329_/A sky130_fd_sc_hd__nand4_4
X_6154_ _7152_/B VGND VGND VPWR VPWR _7042_/C sky130_fd_sc_hd__clkbuf_2
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6085_ _6085_/A _6085_/B VGND VGND VPWR VPWR _6087_/A sky130_fd_sc_hd__xnor2_2
X_5105_ _5105_/A _5105_/B _5104_/X VGND VGND VPWR VPWR _5105_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_85_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5053_/A VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6987_ _6987_/A _6987_/B VGND VGND VPWR VPWR _6988_/C sky130_fd_sc_hd__nand2_1
X_8726_ _8726_/A _8726_/B VGND VGND VPWR VPWR _8727_/B sky130_fd_sc_hd__xnor2_1
XFILLER_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5938_ _5951_/B _5938_/B VGND VGND VPWR VPWR _9056_/A sky130_fd_sc_hd__and2_1
XFILLER_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8657_ _8891_/B VGND VGND VPWR VPWR _9025_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5869_ _7645_/A _6700_/A VGND VGND VPWR VPWR _5871_/A sky130_fd_sc_hd__nand2_1
X_8588_ _8716_/A _9004_/A _8586_/Y _8668_/A VGND VGND VPWR VPWR _8590_/A sky130_fd_sc_hd__o2bb2a_1
X_7608_ _7608_/A _8190_/A VGND VGND VPWR VPWR _7612_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7539_ _7539_/A _7539_/B _7539_/C VGND VGND VPWR VPWR _7539_/Y sky130_fd_sc_hd__nand3_1
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9209_ _9213_/CLK _9209_/D VGND VGND VPWR VPWR _9209_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput67 _9140_/Q VGND VGND VPWR VPWR F[11] sky130_fd_sc_hd__buf_2
Xoutput89 _9160_/Q VGND VGND VPWR VPWR F[31] sky130_fd_sc_hd__buf_2
Xoutput78 _9150_/Q VGND VGND VPWR VPWR F[21] sky130_fd_sc_hd__buf_2
XFILLER_102_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7890_ _7890_/A _7890_/B VGND VGND VPWR VPWR _7891_/C sky130_fd_sc_hd__xnor2_1
X_6910_ _7033_/A _6910_/B VGND VGND VPWR VPWR _6911_/B sky130_fd_sc_hd__xnor2_1
X_6841_ _6740_/C _6845_/B _6838_/Y _6839_/X VGND VGND VPWR VPWR _6843_/C sky130_fd_sc_hd__a211o_1
X_8511_ _8429_/B _8510_/Y _8427_/B VGND VGND VPWR VPWR _8512_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6772_ _6772_/A _6772_/B _6879_/A VGND VGND VPWR VPWR _6940_/B sky130_fd_sc_hd__nor3_4
X_5723_ _9090_/Q _9093_/Q _9088_/Q _4935_/A VGND VGND VPWR VPWR _5723_/X sky130_fd_sc_hd__a22o_1
X_8442_ _8442_/A _8442_/B VGND VGND VPWR VPWR _8444_/B sky130_fd_sc_hd__xnor2_1
X_5654_ _5632_/X _5365_/A _5204_/A _5652_/X _5653_/X VGND VGND VPWR VPWR _9145_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8373_ _8373_/A _8373_/B VGND VGND VPWR VPWR _8492_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4605_ _4605_/A VGND VGND VPWR VPWR _5132_/A sky130_fd_sc_hd__clkbuf_2
X_7324_ _7324_/A _7249_/B VGND VGND VPWR VPWR _7340_/B sky130_fd_sc_hd__or2b_1
X_5585_ _5210_/A _4580_/X _4660_/A _5211_/A _5584_/Y VGND VGND VPWR VPWR _5585_/X
+ sky130_fd_sc_hd__o221a_1
X_4536_ _9109_/Q VGND VGND VPWR VPWR _4737_/A sky130_fd_sc_hd__clkbuf_2
X_7255_ _6775_/A _7852_/C _7252_/Y _7352_/A VGND VGND VPWR VPWR _7256_/B sky130_fd_sc_hd__o2bb2a_1
X_6206_ _6207_/B _6207_/C _6207_/A VGND VGND VPWR VPWR _6210_/A sky130_fd_sc_hd__a21o_1
X_7186_ _7189_/D VGND VGND VPWR VPWR _7186_/Y sky130_fd_sc_hd__clkinv_2
X_6137_ _6760_/A VGND VGND VPWR VPWR _7040_/A sky130_fd_sc_hd__clkbuf_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6068_ _6068_/A _6068_/B _6068_/C VGND VGND VPWR VPWR _6071_/B sky130_fd_sc_hd__nand3_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5019_ _4921_/X _5018_/Y _4799_/A VGND VGND VPWR VPWR _5019_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8709_ _8709_/A _8709_/B VGND VGND VPWR VPWR _8709_/X sky130_fd_sc_hd__or2_1
XFILLER_96_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5370_ _5370_/A _5634_/B VGND VGND VPWR VPWR _5370_/Y sky130_fd_sc_hd__nand2_1
X_7040_ _7040_/A _7153_/D VGND VGND VPWR VPWR _7044_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8991_ _8992_/A _8992_/B VGND VGND VPWR VPWR _9013_/A sky130_fd_sc_hd__or2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7942_ _7942_/A _8046_/B VGND VGND VPWR VPWR _7944_/C sky130_fd_sc_hd__xnor2_1
XFILLER_55_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7873_ _7873_/A _8239_/D VGND VGND VPWR VPWR _7874_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6824_ _9209_/Q VGND VGND VPWR VPWR _7822_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6755_ _7309_/A _6493_/C _7604_/D _7201_/A VGND VGND VPWR VPWR _6756_/B sky130_fd_sc_hd__a22oi_1
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ _5558_/X _4593_/A _5160_/A VGND VGND VPWR VPWR _5706_/Y sky130_fd_sc_hd__a21oi_1
X_8425_ _8328_/B _8336_/X _8423_/Y _8424_/X VGND VGND VPWR VPWR _8510_/B sky130_fd_sc_hd__a211oi_2
X_6686_ _6751_/A _6686_/B VGND VGND VPWR VPWR _6687_/B sky130_fd_sc_hd__xnor2_1
X_5637_ _4661_/A _5389_/X _5368_/X VGND VGND VPWR VPWR _5637_/Y sky130_fd_sc_hd__a21oi_1
X_8356_ _8356_/A _8447_/A VGND VGND VPWR VPWR _8358_/B sky130_fd_sc_hd__or2_1
X_5568_ _5424_/X _4923_/A _5566_/X _5567_/Y _5227_/X VGND VGND VPWR VPWR _5568_/X
+ sky130_fd_sc_hd__a221o_1
X_8287_ _8151_/A _8153_/B _8151_/B VGND VGND VPWR VPWR _8297_/A sky130_fd_sc_hd__o21ba_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7307_ _7307_/A _7307_/B _7822_/C _7307_/D VGND VGND VPWR VPWR _7308_/B sky130_fd_sc_hd__and4_1
X_7238_ _7235_/Y _7319_/A _7237_/X _7160_/B VGND VGND VPWR VPWR _7271_/A sky130_fd_sc_hd__a211o_1
X_5499_ _5315_/A _5403_/X _5497_/X _5498_/Y _5391_/X VGND VGND VPWR VPWR _5499_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7169_ _7170_/A _7281_/C _7167_/X _7168_/Y VGND VGND VPWR VPWR _7171_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4870_ _4960_/B _4869_/X _4870_/S VGND VGND VPWR VPWR _4870_/X sky130_fd_sc_hd__mux2_1
X_6540_ _6585_/A _6585_/B VGND VGND VPWR VPWR _6541_/C sky130_fd_sc_hd__xnor2_1
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6471_ _6377_/A _6377_/B _6376_/B VGND VGND VPWR VPWR _6481_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8210_ _8210_/A _8210_/B VGND VGND VPWR VPWR _8211_/C sky130_fd_sc_hd__nand2_1
X_9190_ _9219_/CLK _9190_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
X_5422_ _5200_/A _5403_/X _5418_/X _5421_/Y _5391_/X VGND VGND VPWR VPWR _5422_/X
+ sky130_fd_sc_hd__a221o_1
X_8141_ _8842_/B VGND VGND VPWR VPWR _8844_/D sky130_fd_sc_hd__buf_2
X_5353_ _5206_/A _5352_/Y _5572_/S VGND VGND VPWR VPWR _5353_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8072_ _8072_/A _8072_/B VGND VGND VPWR VPWR _8076_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5284_ _9069_/Q _5337_/B VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__or2_1
XFILLER_87_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7023_ _7022_/A _7022_/B _7022_/C VGND VGND VPWR VPWR _7161_/A sky130_fd_sc_hd__o21ai_2
XFILLER_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8974_ _8974_/A _9025_/A VGND VGND VPWR VPWR _8974_/Y sky130_fd_sc_hd__nand2_1
X_7925_ _7925_/A VGND VGND VPWR VPWR _8220_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7856_ _7734_/A _7736_/B _7734_/B VGND VGND VPWR VPWR _7857_/B sky130_fd_sc_hd__o21ba_1
X_6807_ _6808_/B _6808_/C _6808_/A VGND VGND VPWR VPWR _6809_/A sky130_fd_sc_hd__a21o_1
X_7787_ _7799_/A _7799_/B VGND VGND VPWR VPWR _7788_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ _5236_/S VGND VGND VPWR VPWR _4999_/X sky130_fd_sc_hd__buf_2
XFILLER_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6738_ _6843_/A _6738_/B VGND VGND VPWR VPWR _6740_/A sky130_fd_sc_hd__nor2_1
X_6669_ _7006_/A _7241_/B _6886_/B _5818_/X VGND VGND VPWR VPWR _6670_/B sky130_fd_sc_hd__a22oi_1
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8408_ _8933_/B VGND VGND VPWR VPWR _8981_/B sky130_fd_sc_hd__buf_2
X_8339_ _8438_/B _8717_/A _8841_/A _8438_/A VGND VGND VPWR VPWR _8343_/A sky130_fd_sc_hd__a22oi_1
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5971_ _5969_/X _5971_/B VGND VGND VPWR VPWR _5974_/A sky130_fd_sc_hd__and2b_1
X_8690_ _8620_/B _8624_/C _8687_/Y _8753_/A VGND VGND VPWR VPWR _8753_/B sky130_fd_sc_hd__a211oi_2
X_7710_ _7710_/A _7818_/B VGND VGND VPWR VPWR _7712_/C sky130_fd_sc_hd__xnor2_1
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4922_ _4767_/A _4960_/B _4963_/B _4921_/X VGND VGND VPWR VPWR _4922_/X sky130_fd_sc_hd__a31o_1
XFILLER_100_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7641_ _8154_/B VGND VGND VPWR VPWR _8721_/B sky130_fd_sc_hd__buf_2
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4853_ _5065_/A _4933_/A VGND VGND VPWR VPWR _4873_/A sky130_fd_sc_hd__nor2_4
X_7572_ _7689_/A _8039_/A _7421_/D _7419_/X VGND VGND VPWR VPWR _7573_/B sky130_fd_sc_hd__a31o_1
X_4784_ _4783_/X _4824_/A _4582_/A VGND VGND VPWR VPWR _4784_/Y sky130_fd_sc_hd__a21oi_1
X_6523_ _6565_/A _6523_/B VGND VGND VPWR VPWR _6524_/B sky130_fd_sc_hd__xnor2_1
X_6454_ _6454_/A _6525_/A VGND VGND VPWR VPWR _6456_/B sky130_fd_sc_hd__xnor2_1
XFILLER_9_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5405_ _5371_/A _9077_/Q _4660_/A _9075_/Q _4572_/A VGND VGND VPWR VPWR _5405_/X
+ sky130_fd_sc_hd__o221a_1
X_9173_ _9218_/CLK input3/X VGND VGND VPWR VPWR _9173_/Q sky130_fd_sc_hd__dfxtp_4
X_6385_ _6385_/A _6385_/B _6480_/B VGND VGND VPWR VPWR _6476_/B sky130_fd_sc_hd__nor3_1
X_8124_ _8125_/A _8125_/B VGND VGND VPWR VPWR _8231_/A sky130_fd_sc_hd__nor2_2
X_5336_ _5287_/X _5335_/X _5336_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
X_8055_ _8056_/A _8056_/B _8056_/C VGND VGND VPWR VPWR _8197_/B sky130_fd_sc_hd__o21a_1
X_5267_ _9081_/Q VGND VGND VPWR VPWR _5604_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7006_ _7006_/A _7006_/B _7348_/B _7119_/C VGND VGND VPWR VPWR _7008_/A sky130_fd_sc_hd__and4_1
XFILLER_75_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5198_ _9067_/Q _5197_/X _5785_/S VGND VGND VPWR VPWR _5199_/A sky130_fd_sc_hd__mux2_1
X_8957_ _8957_/A _8957_/B _8957_/C VGND VGND VPWR VPWR _8958_/B sky130_fd_sc_hd__nor3_1
X_7908_ _8020_/A _8020_/B VGND VGND VPWR VPWR _8022_/A sky130_fd_sc_hd__xnor2_2
X_8888_ _8889_/A _8889_/B VGND VGND VPWR VPWR _8890_/A sky130_fd_sc_hd__nand2_1
X_7839_ _7716_/A _7716_/B _7718_/Y VGND VGND VPWR VPWR _7841_/A sky130_fd_sc_hd__o21bai_1
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6170_ _7347_/A VGND VGND VPWR VPWR _6907_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5121_ _9086_/Q VGND VGND VPWR VPWR _5122_/A sky130_fd_sc_hd__buf_2
X_5052_ _5052_/A _5052_/B VGND VGND VPWR VPWR _5053_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8811_ _8811_/A _8738_/A VGND VGND VPWR VPWR _8812_/A sky130_fd_sc_hd__or2b_1
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8742_ _8742_/A _8812_/B VGND VGND VPWR VPWR _8744_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5954_ _6126_/A _5954_/B _9055_/A VGND VGND VPWR VPWR _9052_/B sky130_fd_sc_hd__nand3_1
X_8673_ _8672_/A _8672_/B _8672_/C VGND VGND VPWR VPWR _8745_/A sky130_fd_sc_hd__a21oi_1
X_4905_ _4905_/A _4905_/B VGND VGND VPWR VPWR _4913_/A sky130_fd_sc_hd__xnor2_4
X_5885_ _5885_/A _5885_/B _5885_/C VGND VGND VPWR VPWR _5896_/B sky130_fd_sc_hd__and3_1
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7624_ _8086_/C VGND VGND VPWR VPWR _8466_/A sky130_fd_sc_hd__clkbuf_2
X_4836_ _4836_/A _4845_/B VGND VGND VPWR VPWR _5074_/A sky130_fd_sc_hd__nor2_1
X_7555_ _8867_/B VGND VGND VPWR VPWR _8909_/B sky130_fd_sc_hd__clkbuf_2
X_6506_ _6563_/B _6506_/B VGND VGND VPWR VPWR _6507_/B sky130_fd_sc_hd__xnor2_2
X_4767_ _4767_/A _4829_/A VGND VGND VPWR VPWR _4787_/B sky130_fd_sc_hd__nor2_4
X_7486_ _7628_/A VGND VGND VPWR VPWR _8069_/A sky130_fd_sc_hd__clkbuf_2
X_4698_ _4864_/A VGND VGND VPWR VPWR _4698_/X sky130_fd_sc_hd__buf_2
X_6437_ _9175_/Q VGND VGND VPWR VPWR _7241_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6368_ _6367_/A _6367_/B _6367_/C VGND VGND VPWR VPWR _6369_/B sky130_fd_sc_hd__o21a_1
X_9156_ _9218_/CLK _9156_/D VGND VGND VPWR VPWR _9156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8107_ _8107_/A _8107_/B VGND VGND VPWR VPWR _8135_/A sky130_fd_sc_hd__and2_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5319_ _4585_/A _5404_/A _5219_/X VGND VGND VPWR VPWR _5319_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_88_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6299_ _6304_/A _6304_/B _6304_/C VGND VGND VPWR VPWR _6300_/B sky130_fd_sc_hd__a21oi_1
X_9087_ _9090_/CLK _9087_/D VGND VGND VPWR VPWR _9087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8038_ _8038_/A VGND VGND VPWR VPWR _8322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 _9143_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _4560_/A _5669_/X _5670_/S VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4621_ _4541_/X _4617_/X _5765_/C VGND VGND VPWR VPWR _4621_/X sky130_fd_sc_hd__o21a_1
X_7340_ _7340_/A _7340_/B _7340_/C VGND VGND VPWR VPWR _7340_/X sky130_fd_sc_hd__and3_1
X_4552_ _9102_/Q VGND VGND VPWR VPWR _5733_/S sky130_fd_sc_hd__clkinv_2
X_7271_ _7271_/A _7319_/B _7271_/C _7383_/A VGND VGND VPWR VPWR _7383_/B sky130_fd_sc_hd__nand4_1
XFILLER_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9010_ _9009_/A _9009_/B _9009_/C VGND VGND VPWR VPWR _9011_/B sky130_fd_sc_hd__a21oi_1
X_6222_ _6213_/Y _6304_/A VGND VGND VPWR VPWR _6385_/A sky130_fd_sc_hd__nand2b_1
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6153_ _9172_/Q VGND VGND VPWR VPWR _7152_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _7569_/C _7499_/A VGND VGND VPWR VPWR _6085_/B sky130_fd_sc_hd__nand2_1
X_5104_ _4972_/Y _5019_/X _5067_/X _5391_/A VGND VGND VPWR VPWR _5104_/X sky130_fd_sc_hd__a31o_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5035_ _5035_/A _5035_/B VGND VGND VPWR VPWR _5053_/A sky130_fd_sc_hd__nor2_2
XFILLER_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6986_ _6986_/A _6986_/B _6986_/C VGND VGND VPWR VPWR _6987_/B sky130_fd_sc_hd__nand3_1
X_8725_ _8725_/A _8787_/B VGND VGND VPWR VPWR _8726_/B sky130_fd_sc_hd__nor2_1
X_5937_ _5897_/A _5896_/B _9060_/A VGND VGND VPWR VPWR _5938_/B sky130_fd_sc_hd__o21bai_1
X_8656_ _8656_/A _8641_/B VGND VGND VPWR VPWR _8705_/B sky130_fd_sc_hd__or2b_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7607_ _7728_/C VGND VGND VPWR VPWR _8190_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5868_ _6361_/B VGND VGND VPWR VPWR _6700_/A sky130_fd_sc_hd__buf_2
X_8587_ _8587_/A _8587_/B _8660_/C VGND VGND VPWR VPWR _8668_/A sky130_fd_sc_hd__and3_1
X_5799_ _9165_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__clkbuf_2
X_4819_ _4928_/A VGND VGND VPWR VPWR _4914_/A sky130_fd_sc_hd__inv_2
X_7538_ _7538_/A _7668_/A _7536_/Y VGND VGND VPWR VPWR _7668_/B sky130_fd_sc_hd__nor3b_2
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7469_ _7469_/A _7469_/B VGND VGND VPWR VPWR _7470_/B sky130_fd_sc_hd__nor2_1
X_9208_ _9208_/CLK _9208_/D VGND VGND VPWR VPWR _9208_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput79 _9151_/Q VGND VGND VPWR VPWR F[22] sky130_fd_sc_hd__buf_2
Xoutput68 _9141_/Q VGND VGND VPWR VPWR F[12] sky130_fd_sc_hd__buf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9139_ _9220_/CLK _9139_/D VGND VGND VPWR VPWR _9139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6840_ _6838_/Y _6839_/X _6740_/C _6845_/B VGND VGND VPWR VPWR _6843_/B sky130_fd_sc_hd__o211ai_2
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ _6772_/B _6879_/A _6772_/A VGND VGND VPWR VPWR _6940_/A sky130_fd_sc_hd__o21a_1
XFILLER_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8510_ _8510_/A _8510_/B VGND VGND VPWR VPWR _8510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5722_ _5765_/C _5365_/A _5278_/X _4812_/X _5721_/X VGND VGND VPWR VPWR _9148_/D
+ sky130_fd_sc_hd__o221ai_1
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8441_ _8584_/A _8792_/A VGND VGND VPWR VPWR _8442_/B sky130_fd_sc_hd__nand2_1
X_5653_ _5653_/A _5653_/B VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__or2_1
X_8372_ _8568_/A _8846_/B VGND VGND VPWR VPWR _8373_/B sky130_fd_sc_hd__nand2_1
X_5584_ _5144_/A _5607_/A _4847_/A VGND VGND VPWR VPWR _5584_/Y sky130_fd_sc_hd__a21oi_1
X_4604_ _4774_/A VGND VGND VPWR VPWR _4605_/A sky130_fd_sc_hd__clkbuf_2
X_4535_ _4535_/A VGND VGND VPWR VPWR _4535_/X sky130_fd_sc_hd__clkbuf_2
X_7323_ _7209_/B _7321_/X _7319_/X _7533_/A VGND VGND VPWR VPWR _7533_/B sky130_fd_sc_hd__a211oi_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7254_ _7252_/Y _7352_/A _7254_/C _7254_/D VGND VGND VPWR VPWR _7352_/B sky130_fd_sc_hd__and4bb_1
XFILLER_104_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6205_ _6292_/A _6205_/B VGND VGND VPWR VPWR _6207_/A sky130_fd_sc_hd__nor2_1
X_7185_ _6251_/A _7419_/C _7419_/D _6361_/B VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__a22o_1
X_6136_ _9170_/Q VGND VGND VPWR VPWR _6760_/A sky130_fd_sc_hd__clkbuf_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6068_/B _6068_/C _6068_/A VGND VGND VPWR VPWR _6071_/A sky130_fd_sc_hd__a21o_1
XFILLER_73_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5018_ _5177_/A _4964_/X _5017_/Y _4967_/X VGND VGND VPWR VPWR _5018_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6969_ _7099_/A VGND VGND VPWR VPWR _6986_/B sky130_fd_sc_hd__inv_2
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8708_ _8637_/B _8640_/B _8705_/X _8768_/A VGND VGND VPWR VPWR _8768_/B sky130_fd_sc_hd__a211oi_2
X_8639_ _8639_/A _8639_/B _8639_/C VGND VGND VPWR VPWR _8640_/B sky130_fd_sc_hd__nand3_1
XFILLER_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8990_ _8990_/A _8990_/B VGND VGND VPWR VPWR _8992_/B sky130_fd_sc_hd__xor2_1
XFILLER_82_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7941_ _8047_/C _7941_/B VGND VGND VPWR VPWR _8046_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7872_ _7966_/D VGND VGND VPWR VPWR _8239_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6823_ _9208_/Q VGND VGND VPWR VPWR _6825_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6754_ _7419_/A _6754_/B _7728_/B _7222_/D VGND VGND VPWR VPWR _6756_/A sky130_fd_sc_hd__and4_1
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6685_ _6751_/B _6805_/B VGND VGND VPWR VPWR _6686_/B sky130_fd_sc_hd__nor2_1
X_5705_ _5287_/A _5154_/X _5704_/X _5249_/A VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__a211o_1
X_8424_ _8423_/A _8423_/B _8423_/C VGND VGND VPWR VPWR _8424_/X sky130_fd_sc_hd__o21a_1
X_5636_ _4650_/A _5205_/A _5634_/Y _5635_/X _4661_/A VGND VGND VPWR VPWR _5636_/X
+ sky130_fd_sc_hd__a221o_1
X_8355_ _8355_/A _8355_/B VGND VGND VPWR VPWR _8447_/A sky130_fd_sc_hd__and2_1
X_5567_ _5393_/A _4556_/A _5213_/A VGND VGND VPWR VPWR _5567_/Y sky130_fd_sc_hd__a21oi_1
X_8286_ _8286_/A _8286_/B VGND VGND VPWR VPWR _8307_/A sky130_fd_sc_hd__xor2_1
X_7306_ _6925_/A _6825_/C _7706_/D _7037_/A VGND VGND VPWR VPWR _7308_/A sky130_fd_sc_hd__a22oi_1
X_5498_ _5450_/X _5126_/X _5181_/X VGND VGND VPWR VPWR _5498_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7237_ _7157_/B _7237_/B VGND VGND VPWR VPWR _7237_/X sky130_fd_sc_hd__and2b_1
XFILLER_77_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7168_ _7053_/C _7053_/Y _7165_/Y _7274_/B VGND VGND VPWR VPWR _7168_/Y sky130_fd_sc_hd__o211ai_2
X_6119_ _6119_/A _6119_/B VGND VGND VPWR VPWR _6213_/A sky130_fd_sc_hd__nor2_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7099_ _7099_/A _7099_/B VGND VGND VPWR VPWR _7100_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6470_ _6470_/A _6470_/B VGND VGND VPWR VPWR _6481_/A sky130_fd_sc_hd__xnor2_2
X_5421_ _5271_/X _5420_/X _4629_/A VGND VGND VPWR VPWR _5421_/Y sky130_fd_sc_hd__a21oi_1
X_8140_ _8664_/D VGND VGND VPWR VPWR _8842_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5352_ _4726_/X _5278_/X _5351_/X VGND VGND VPWR VPWR _5352_/Y sky130_fd_sc_hd__o21ai_1
X_8071_ _8071_/A _8349_/B _8071_/C VGND VGND VPWR VPWR _8072_/B sky130_fd_sc_hd__and3_1
XFILLER_99_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7022_ _7022_/A _7022_/B _7022_/C VGND VGND VPWR VPWR _7024_/A sky130_fd_sc_hd__or3_1
X_5283_ _5200_/X _5282_/X _5336_/S VGND VGND VPWR VPWR _5283_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8973_ _8961_/A _8973_/B VGND VGND VPWR VPWR _8973_/X sky130_fd_sc_hd__and2b_1
X_7924_ _7924_/A _7924_/B VGND VGND VPWR VPWR _7927_/A sky130_fd_sc_hd__nor2_1
X_7855_ _7855_/A _7855_/B VGND VGND VPWR VPWR _7978_/B sky130_fd_sc_hd__xnor2_1
X_6806_ _6934_/B _6806_/B VGND VGND VPWR VPWR _6808_/A sky130_fd_sc_hd__and2_1
X_7786_ _7786_/A _7903_/A VGND VGND VPWR VPWR _7799_/B sky130_fd_sc_hd__and2_1
X_4998_ _4998_/A VGND VGND VPWR VPWR _5028_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6737_ _6737_/A _6737_/B _6737_/C VGND VGND VPWR VPWR _6738_/B sky130_fd_sc_hd__and3_1
X_6668_ _6894_/A _7119_/B _7131_/C _7131_/D VGND VGND VPWR VPWR _6670_/A sky130_fd_sc_hd__and4_1
X_8407_ _8267_/B _8405_/X _8490_/B _8404_/Y VGND VGND VPWR VPWR _8419_/B sky130_fd_sc_hd__a211oi_4
X_6599_ _6599_/A _6658_/A VGND VGND VPWR VPWR _6659_/B sky130_fd_sc_hd__xnor2_1
X_5619_ _5618_/X _5129_/X _5175_/X VGND VGND VPWR VPWR _5619_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8338_ _8607_/D VGND VGND VPWR VPWR _8841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8269_ _8269_/A VGND VGND VPWR VPWR _8792_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5970_ _9165_/Q _6885_/A _9169_/Q _6235_/A VGND VGND VPWR VPWR _5971_/B sky130_fd_sc_hd__a22o_1
X_4921_ _4844_/X _4971_/B _4834_/A VGND VGND VPWR VPWR _4921_/X sky130_fd_sc_hd__a21o_1
X_7640_ _7640_/A VGND VGND VPWR VPWR _8154_/B sky130_fd_sc_hd__clkbuf_2
X_4852_ _4852_/A _4852_/B VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__and2_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7571_ _7571_/A VGND VGND VPWR VPWR _8039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4783_ _4783_/A VGND VGND VPWR VPWR _4783_/X sky130_fd_sc_hd__buf_2
X_6522_ _6565_/B _6611_/B VGND VGND VPWR VPWR _6523_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6453_ _6328_/A _6327_/B _6327_/A VGND VGND VPWR VPWR _6525_/A sky130_fd_sc_hd__o21ba_1
X_9172_ _9212_/CLK input2/X VGND VGND VPWR VPWR _9172_/Q sky130_fd_sc_hd__dfxtp_1
X_5404_ _5404_/A _5634_/B VGND VGND VPWR VPWR _5404_/Y sky130_fd_sc_hd__nand2_1
X_8123_ _8016_/A _8016_/B _8122_/X VGND VGND VPWR VPWR _8125_/B sky130_fd_sc_hd__a21boi_1
X_6384_ _6302_/A _6302_/B _6304_/Y _6300_/B _6383_/B VGND VGND VPWR VPWR _6476_/A
+ sky130_fd_sc_hd__a311oi_2
X_5335_ _5245_/X _5334_/X _5428_/S VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__mux2_1
X_8054_ _8054_/A _8184_/B VGND VGND VPWR VPWR _8056_/C sky130_fd_sc_hd__xnor2_1
X_5266_ _5414_/A VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7005_ _7118_/A _8091_/C VGND VGND VPWR VPWR _7009_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5197_ _5510_/A _5117_/X _5196_/X VGND VGND VPWR VPWR _5197_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8956_ _8957_/A _8957_/B _8957_/C VGND VGND VPWR VPWR _8958_/A sky130_fd_sc_hd__o21a_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7907_ _7791_/A _7791_/B _7790_/B VGND VGND VPWR VPWR _8020_/B sky130_fd_sc_hd__a21oi_2
X_8887_ _8887_/A _8937_/B VGND VGND VPWR VPWR _8889_/B sky130_fd_sc_hd__or2_1
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7838_ _7915_/A VGND VGND VPWR VPWR _7841_/C sky130_fd_sc_hd__inv_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7769_ _7769_/A VGND VGND VPWR VPWR _8349_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_105_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5120_ _5120_/A VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__buf_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5051_ _5053_/A _5051_/B VGND VGND VPWR VPWR _5051_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8810_ _8810_/A _8872_/A VGND VGND VPWR VPWR _8830_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8741_ _8741_/A _8741_/B VGND VGND VPWR VPWR _8812_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ _9057_/A _9054_/B VGND VGND VPWR VPWR _9055_/A sky130_fd_sc_hd__nor2_1
X_8672_ _8672_/A _8672_/B _8672_/C VGND VGND VPWR VPWR _8686_/B sky130_fd_sc_hd__and3_1
X_4904_ _4991_/A _4904_/B VGND VGND VPWR VPWR _4905_/B sky130_fd_sc_hd__nand2_1
X_5884_ _5885_/B _5885_/C _5885_/A VGND VGND VPWR VPWR _5897_/A sky130_fd_sc_hd__a21oi_2
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7623_ _7873_/A VGND VGND VPWR VPWR _8137_/A sky130_fd_sc_hd__clkbuf_2
X_4835_ _4929_/A _4914_/A VGND VGND VPWR VPWR _4927_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7554_ _7071_/A _7071_/B _7071_/C _7552_/Y _7553_/X VGND VGND VPWR VPWR _7677_/C
+ sky130_fd_sc_hd__a311o_2
X_4766_ _4842_/A _4824_/A VGND VGND VPWR VPWR _4829_/A sky130_fd_sc_hd__and2_1
X_6505_ _6407_/A _6406_/A _6406_/B VGND VGND VPWR VPWR _6506_/B sky130_fd_sc_hd__o21ba_1
X_7485_ _7485_/A _8086_/C VGND VGND VPWR VPWR _7492_/A sky130_fd_sc_hd__nand2_1
X_4697_ _4697_/A VGND VGND VPWR VPWR _4889_/A sky130_fd_sc_hd__clkbuf_2
X_6436_ _7153_/C VGND VGND VPWR VPWR _7583_/B sky130_fd_sc_hd__clkbuf_2
X_9224_ _9224_/CLK hold14/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
X_9155_ _9220_/CLK _9155_/D VGND VGND VPWR VPWR _9155_/Q sky130_fd_sc_hd__dfxtp_1
X_6367_ _6367_/A _6367_/B _6367_/C VGND VGND VPWR VPWR _6369_/A sky130_fd_sc_hd__nor3_1
X_8106_ _8105_/B _8203_/B _8105_/A VGND VGND VPWR VPWR _8107_/B sky130_fd_sc_hd__a21o_1
X_5318_ _4847_/A _9075_/Q _5316_/Y _5317_/X _4584_/A VGND VGND VPWR VPWR _5318_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6298_ _6304_/A _6304_/B _6304_/C VGND VGND VPWR VPWR _6300_/A sky130_fd_sc_hd__and3_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_9086_ _9090_/CLK _9086_/D VGND VGND VPWR VPWR _9086_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8037_ _8037_/A _8037_/B VGND VGND VPWR VPWR _8041_/A sky130_fd_sc_hd__nor2_1
X_5249_ _5249_/A VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8939_ _8985_/A _8939_/B VGND VGND VPWR VPWR _8942_/B sky130_fd_sc_hd__or2_1
XFILLER_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _5695_/S VGND VGND VPWR VPWR _5765_/C sky130_fd_sc_hd__clkbuf_2
X_4551_ _4608_/B VGND VGND VPWR VPWR _5754_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7270_ _7139_/C _7140_/B _7267_/X _7268_/Y VGND VGND VPWR VPWR _7383_/A sky130_fd_sc_hd__a211o_2
X_6221_ _6221_/A _6221_/B VGND VGND VPWR VPWR _6304_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6152_ _6702_/A VGND VGND VPWR VPWR _6922_/B sky130_fd_sc_hd__clkbuf_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5103_/A VGND VGND VPWR VPWR _5105_/A sky130_fd_sc_hd__buf_2
XFILLER_97_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6083_ _6660_/A VGND VGND VPWR VPWR _7499_/A sky130_fd_sc_hd__buf_2
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5033_/A _5033_/B _5033_/C VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__o21a_1
XFILLER_38_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6985_ _6986_/A _6986_/B _6986_/C VGND VGND VPWR VPWR _6987_/A sky130_fd_sc_hd__a21o_1
X_8724_ _8724_/A _8841_/A _8724_/C VGND VGND VPWR VPWR _8787_/B sky130_fd_sc_hd__and3_1
X_5936_ _5952_/A _5951_/B _5933_/X _6047_/A VGND VGND VPWR VPWR _5954_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8655_ _8655_/A VGND VGND VPWR VPWR _9101_/D sky130_fd_sc_hd__clkbuf_1
X_7606_ _7606_/A _7606_/B VGND VGND VPWR VPWR _7615_/A sky130_fd_sc_hd__xnor2_2
X_5867_ _6593_/A VGND VGND VPWR VPWR _7645_/A sky130_fd_sc_hd__buf_4
X_8586_ _8438_/A _8780_/B _8660_/C VGND VGND VPWR VPWR _8586_/Y sky130_fd_sc_hd__a21oi_1
X_4818_ _4852_/B VGND VGND VPWR VPWR _4928_/A sky130_fd_sc_hd__clkbuf_2
X_5798_ _7201_/A _5945_/A _7766_/A _5922_/A VGND VGND VPWR VPWR _5898_/C sky130_fd_sc_hd__and4_2
X_4749_ _9123_/Q _9115_/Q VGND VGND VPWR VPWR _4750_/B sky130_fd_sc_hd__or2_1
X_7537_ _7538_/A _7668_/A _7536_/Y VGND VGND VPWR VPWR _7537_/X sky130_fd_sc_hd__o21ba_1
X_7468_ _8091_/A _8243_/A _8050_/B _7847_/D VGND VGND VPWR VPWR _7469_/B sky130_fd_sc_hd__and4_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9207_ _9220_/CLK _9207_/D VGND VGND VPWR VPWR _9207_/Q sky130_fd_sc_hd__dfxtp_2
X_6419_ _6414_/X _6417_/X _6411_/X _6413_/Y VGND VGND VPWR VPWR _6483_/C sky130_fd_sc_hd__o211a_1
X_7399_ _7539_/A _7539_/B _7539_/C VGND VGND VPWR VPWR _7399_/X sky130_fd_sc_hd__and3_1
Xoutput69 _9142_/Q VGND VGND VPWR VPWR F[13] sky130_fd_sc_hd__buf_2
XFILLER_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9138_ _9199_/CLK _9138_/D VGND VGND VPWR VPWR _9138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9069_ _9090_/CLK _9069_/D VGND VGND VPWR VPWR _9069_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6770_ _6709_/A _6709_/B _6769_/X VGND VGND VPWR VPWR _6772_/A sky130_fd_sc_hd__a21oi_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5721_ _4999_/X _4535_/X _5719_/X _5720_/Y _5511_/A VGND VGND VPWR VPWR _5721_/X
+ sky130_fd_sc_hd__a221o_1
X_8440_ _8717_/A VGND VGND VPWR VPWR _8792_/A sky130_fd_sc_hd__clkbuf_2
X_5652_ _5606_/X _5651_/X _5698_/S VGND VGND VPWR VPWR _5652_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8371_ _8371_/A VGND VGND VPWR VPWR _8568_/A sky130_fd_sc_hd__clkbuf_2
X_5583_ _5754_/A VGND VGND VPWR VPWR _5583_/X sky130_fd_sc_hd__clkbuf_2
X_4603_ _9101_/Q VGND VGND VPWR VPWR _4774_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7322_ _7319_/X _7533_/A _7209_/B _7321_/X VGND VGND VPWR VPWR _7386_/A sky130_fd_sc_hd__o211a_1
X_4534_ _9111_/Q VGND VGND VPWR VPWR _4535_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7253_ _7253_/A _7253_/B _9179_/Q _9183_/Q VGND VGND VPWR VPWR _7352_/A sky130_fd_sc_hd__and4_1
X_7184_ _9213_/Q VGND VGND VPWR VPWR _7571_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6204_ _6204_/A _6204_/B _6204_/C VGND VGND VPWR VPWR _6205_/B sky130_fd_sc_hd__and3_1
X_6135_ _7307_/B VGND VGND VPWR VPWR _6607_/A sky130_fd_sc_hd__buf_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6066_ _7257_/A _7148_/B VGND VGND VPWR VPWR _6068_/A sky130_fd_sc_hd__and2_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5017_ _5385_/A _5017_/B VGND VGND VPWR VPWR _5017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8707_ _8705_/X _8768_/A _8637_/B _8640_/B VGND VGND VPWR VPWR _8707_/X sky130_fd_sc_hd__o211a_1
X_6968_ _6968_/A _6968_/B _7923_/C _8175_/D VGND VGND VPWR VPWR _7099_/A sky130_fd_sc_hd__and4_1
X_6899_ _6899_/A _6993_/A VGND VGND VPWR VPWR _6994_/B sky130_fd_sc_hd__xnor2_1
X_5919_ _9198_/Q VGND VGND VPWR VPWR _7361_/C sky130_fd_sc_hd__clkbuf_4
X_8638_ _8639_/A _8756_/B _8639_/C VGND VGND VPWR VPWR _8640_/A sky130_fd_sc_hd__a21o_1
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8569_ _8569_/A _8569_/B VGND VGND VPWR VPWR _8571_/C sky130_fd_sc_hd__xor2_1
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7940_ _8036_/B _7940_/B VGND VGND VPWR VPWR _7941_/B sky130_fd_sc_hd__nand2_1
X_7871_ _7754_/B _8068_/A _7870_/X VGND VGND VPWR VPWR _7874_/A sky130_fd_sc_hd__a21oi_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6822_ _7187_/B _7938_/C VGND VGND VPWR VPWR _6822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6753_ _7187_/A _7730_/B VGND VGND VPWR VPWR _6757_/A sky130_fd_sc_hd__nand2_1
X_6684_ _7808_/B _7988_/A _6684_/C VGND VGND VPWR VPWR _6805_/B sky130_fd_sc_hd__and3_1
X_5704_ _9091_/Q _5618_/A _5702_/Y _5703_/X _4566_/A VGND VGND VPWR VPWR _5704_/X
+ sky130_fd_sc_hd__o221a_1
X_8423_ _8423_/A _8423_/B _8423_/C VGND VGND VPWR VPWR _8423_/Y sky130_fd_sc_hd__nor3_1
X_5635_ _5558_/A _5122_/A _4676_/C _5124_/A _4572_/A VGND VGND VPWR VPWR _5635_/X
+ sky130_fd_sc_hd__o221a_1
X_8354_ _8355_/A _8355_/B VGND VGND VPWR VPWR _8356_/A sky130_fd_sc_hd__nor2_1
X_5566_ _5214_/X _5420_/A _5564_/X _5565_/Y _5001_/A VGND VGND VPWR VPWR _5566_/X
+ sky130_fd_sc_hd__a221o_1
X_8285_ _8415_/A _8898_/B VGND VGND VPWR VPWR _8286_/B sky130_fd_sc_hd__nand2_1
X_7305_ _7224_/A _7223_/A _7223_/B VGND VGND VPWR VPWR _7311_/A sky130_fd_sc_hd__o21ba_1
X_5497_ _5245_/A _5177_/X _5495_/X _5496_/Y _5126_/A VGND VGND VPWR VPWR _5497_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7236_ _7235_/A _7235_/B _7235_/C VGND VGND VPWR VPWR _7319_/A sky130_fd_sc_hd__a21o_2
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7167_ _7165_/Y _7274_/B _7053_/C _7053_/Y VGND VGND VPWR VPWR _7167_/X sky130_fd_sc_hd__a211o_1
XFILLER_100_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6118_ _6118_/A _6118_/B _6118_/C VGND VGND VPWR VPWR _6119_/B sky130_fd_sc_hd__and3_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7099_/A _7099_/B VGND VGND VPWR VPWR _7281_/A sky130_fd_sc_hd__and2_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6049_ _9052_/A _9052_/C _6049_/C _6125_/A VGND VGND VPWR VPWR _6051_/A sky130_fd_sc_hd__and4bb_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5420_ _5420_/A VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__buf_2
X_5351_ _4721_/X _5189_/X _5349_/X _5350_/Y _5230_/X VGND VGND VPWR VPWR _5351_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8070_ _8071_/A _8587_/B _8071_/C VGND VGND VPWR VPWR _8072_/A sky130_fd_sc_hd__a21oi_1
X_5282_ _5117_/X _5281_/X _5282_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
X_7021_ _7021_/A _7021_/B VGND VGND VPWR VPWR _7022_/C sky130_fd_sc_hd__xnor2_1
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8972_ _8972_/A _8972_/B VGND VGND VPWR VPWR _9107_/D sky130_fd_sc_hd__xor2_1
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7923_ _8038_/A _7923_/B _7923_/C _7923_/D VGND VGND VPWR VPWR _7924_/B sky130_fd_sc_hd__and4_1
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7854_ _8093_/A _8086_/C VGND VGND VPWR VPWR _7855_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7785_ _7784_/A _7784_/B _7784_/C VGND VGND VPWR VPWR _7903_/A sky130_fd_sc_hd__o21ai_1
X_6805_ _6805_/A _6805_/B _6805_/C VGND VGND VPWR VPWR _6806_/B sky130_fd_sc_hd__or3_1
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6736_ _6737_/A _6737_/B _6737_/C VGND VGND VPWR VPWR _6843_/A sky130_fd_sc_hd__a21oi_2
X_4997_ _5067_/A VGND VGND VPWR VPWR _4998_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6667_ _6667_/A VGND VGND VPWR VPWR _7119_/B sky130_fd_sc_hd__buf_2
X_8406_ _8490_/B _8404_/Y _8267_/B _8405_/X VGND VGND VPWR VPWR _8419_/A sky130_fd_sc_hd__o211a_1
X_6598_ _6537_/A _6536_/B _6536_/A VGND VGND VPWR VPWR _6658_/A sky130_fd_sc_hd__o21ba_1
X_5618_ _5618_/A VGND VGND VPWR VPWR _5618_/X sky130_fd_sc_hd__clkbuf_4
X_8337_ _8337_/A VGND VGND VPWR VPWR _8438_/B sky130_fd_sc_hd__clkbuf_2
X_5549_ _5364_/A _5403_/X _5547_/X _5548_/Y _5391_/X VGND VGND VPWR VPWR _5549_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8268_ _8268_/A VGND VGND VPWR VPWR _8452_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8199_ _8199_/A _8199_/B VGND VGND VPWR VPWR _8201_/B sky130_fd_sc_hd__nand2_1
X_7219_ _7219_/A _7137_/B VGND VGND VPWR VPWR _7235_/B sky130_fd_sc_hd__or2b_1
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _4920_/A VGND VGND VPWR VPWR _4963_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4851_ _4852_/A _4928_/A VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__nor2_2
X_7570_ _7570_/A _7570_/B VGND VGND VPWR VPWR _7573_/A sky130_fd_sc_hd__nor2_1
X_4782_ _5656_/B _4769_/B _4781_/X VGND VGND VPWR VPWR _4782_/X sky130_fd_sc_hd__a21o_1
X_6521_ _7694_/A _7988_/A _6521_/C VGND VGND VPWR VPWR _6611_/B sky130_fd_sc_hd__and3_1
XFILLER_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6452_ _6452_/A _6452_/B VGND VGND VPWR VPWR _6454_/A sky130_fd_sc_hd__xnor2_2
X_9171_ _9213_/CLK _9171_/D VGND VGND VPWR VPWR _9171_/Q sky130_fd_sc_hd__dfxtp_2
X_5403_ _5403_/A VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8122_ _8122_/A _8015_/B VGND VGND VPWR VPWR _8122_/X sky130_fd_sc_hd__or2b_1
X_6383_ _6383_/A _6383_/B VGND VGND VPWR VPWR _9079_/D sky130_fd_sc_hd__xnor2_1
X_5334_ _5200_/X _5333_/X _5427_/S VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__mux2_1
X_8053_ _8053_/A _8053_/B VGND VGND VPWR VPWR _8184_/B sky130_fd_sc_hd__xnor2_1
X_5265_ _5132_/X _5246_/Y _5262_/X _5264_/Y _4642_/A VGND VGND VPWR VPWR _5265_/X
+ sky130_fd_sc_hd__a221o_1
X_7004_ _7119_/D VGND VGND VPWR VPWR _8091_/C sky130_fd_sc_hd__buf_2
X_5196_ _4535_/A _5120_/X _5191_/X _5195_/Y _9112_/Q VGND VGND VPWR VPWR _5196_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8955_ _8955_/A _8955_/B VGND VGND VPWR VPWR _8957_/C sky130_fd_sc_hd__nand2_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7906_ _7911_/A _7911_/B VGND VGND VPWR VPWR _8020_/A sky130_fd_sc_hd__xnor2_2
X_8886_ _8886_/A VGND VGND VPWR VPWR _9105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7837_ _7837_/A _7837_/B _7837_/C VGND VGND VPWR VPWR _7915_/A sky130_fd_sc_hd__and3_1
XFILLER_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7768_ _7984_/A _7643_/B _7876_/A VGND VGND VPWR VPWR _7771_/A sky130_fd_sc_hd__a21o_1
X_7699_ _7699_/A _7699_/B VGND VGND VPWR VPWR _7702_/A sky130_fd_sc_hd__xor2_1
X_6719_ _6719_/A _6719_/B VGND VGND VPWR VPWR _6737_/B sky130_fd_sc_hd__or2_1
XFILLER_3_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5050_ _5052_/B _5050_/B VGND VGND VPWR VPWR _5051_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8740_ _8741_/A _8741_/B VGND VGND VPWR VPWR _8742_/A sky130_fd_sc_hd__or2_1
X_5952_ _5952_/A _5952_/B VGND VGND VPWR VPWR _9054_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4903_ _9125_/Q _9117_/Q VGND VGND VPWR VPWR _4904_/B sky130_fd_sc_hd__or2_1
X_8671_ _8671_/A _8671_/B VGND VGND VPWR VPWR _8672_/C sky130_fd_sc_hd__xnor2_1
X_5883_ _5883_/A _5883_/B VGND VGND VPWR VPWR _5885_/A sky130_fd_sc_hd__xnor2_1
X_7622_ _7622_/A _7622_/B VGND VGND VPWR VPWR _7660_/A sky130_fd_sc_hd__and2_1
X_4834_ _4834_/A VGND VGND VPWR VPWR _5714_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7553_ _7553_/A _7553_/B _7408_/A VGND VGND VPWR VPWR _7553_/X sky130_fd_sc_hd__or3b_1
X_4765_ _4842_/A _4842_/B VGND VGND VPWR VPWR _4767_/A sky130_fd_sc_hd__nor2_1
X_6504_ _6504_/A _6504_/B VGND VGND VPWR VPWR _6563_/B sky130_fd_sc_hd__xnor2_2
X_7484_ _7959_/D VGND VGND VPWR VPWR _8086_/C sky130_fd_sc_hd__buf_2
X_9223_ _9223_/CLK _9223_/D VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
X_4696_ _5103_/A VGND VGND VPWR VPWR _4697_/A sky130_fd_sc_hd__clkbuf_2
X_6435_ _7499_/A _7808_/B VGND VGND VPWR VPWR _6445_/A sky130_fd_sc_hd__nand2_1
X_9154_ _9210_/CLK _9154_/D VGND VGND VPWR VPWR _9154_/Q sky130_fd_sc_hd__dfxtp_1
X_6366_ _6366_/A _6417_/C VGND VGND VPWR VPWR _6367_/C sky130_fd_sc_hd__xnor2_1
X_8105_ _8105_/A _8105_/B _8203_/B VGND VGND VPWR VPWR _8107_/A sky130_fd_sc_hd__nand3_1
X_5317_ _5252_/A _9074_/Q _4659_/A _9072_/Q _4706_/S VGND VGND VPWR VPWR _5317_/X
+ sky130_fd_sc_hd__o221a_1
X_9085_ _9090_/CLK _9085_/D VGND VGND VPWR VPWR _9085_/Q sky130_fd_sc_hd__dfxtp_1
X_8036_ _8177_/A _8036_/B _8269_/A _8175_/D VGND VGND VPWR VPWR _8037_/B sky130_fd_sc_hd__and4_1
X_6297_ _6385_/A _6385_/B VGND VGND VPWR VPWR _6304_/C sky130_fd_sc_hd__xor2_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5248_ _5248_/A VGND VGND VPWR VPWR _5248_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5179_ _5179_/A VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__buf_2
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8938_ _8937_/A _8937_/B _8937_/C VGND VGND VPWR VPWR _8939_/B sky130_fd_sc_hd__o21a_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8869_ _8870_/A _8870_/B VGND VGND VPWR VPWR _8913_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _4550_/A VGND VGND VPWR VPWR _4608_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6220_ _6220_/A VGND VGND VPWR VPWR _9077_/D sky130_fd_sc_hd__clkbuf_1
X_6151_ _6151_/A _6572_/B _6778_/B _7706_/B VGND VGND VPWR VPWR _6157_/A sky130_fd_sc_hd__and4_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A VGND VGND VPWR VPWR _9158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _7293_/B VGND VGND VPWR VPWR _7569_/C sky130_fd_sc_hd__clkbuf_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B _5033_/C VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__nor3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6984_ _7106_/A _6984_/B VGND VGND VPWR VPWR _6986_/C sky130_fd_sc_hd__xnor2_1
X_8723_ _8666_/A _8844_/B _8724_/C VGND VGND VPWR VPWR _8725_/A sky130_fd_sc_hd__a21oi_1
X_5935_ _5952_/A _5951_/B _5933_/X _6047_/A VGND VGND VPWR VPWR _6126_/A sky130_fd_sc_hd__or4bb_1
X_5866_ _7365_/A VGND VGND VPWR VPWR _6593_/A sky130_fd_sc_hd__clkbuf_2
X_8654_ _8652_/X _8714_/B VGND VGND VPWR VPWR _8655_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7605_ _7605_/A _7605_/B VGND VGND VPWR VPWR _7606_/B sky130_fd_sc_hd__nor2_1
X_4817_ _4816_/B _4828_/C _4817_/S VGND VGND VPWR VPWR _4852_/B sky130_fd_sc_hd__mux2_1
X_8585_ _8844_/D VGND VGND VPWR VPWR _9004_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5797_ _9162_/Q VGND VGND VPWR VPWR _5922_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4748_ _9123_/Q _9115_/Q VGND VGND VPWR VPWR _4816_/A sky130_fd_sc_hd__nand2_2
X_7536_ _7536_/A _7536_/B VGND VGND VPWR VPWR _7536_/Y sky130_fd_sc_hd__xnor2_1
X_7467_ _8091_/B _8050_/B _8190_/B _8154_/A VGND VGND VPWR VPWR _7469_/A sky130_fd_sc_hd__a22oi_1
X_4679_ _4535_/X _4625_/X _5511_/A VGND VGND VPWR VPWR _4680_/B sky130_fd_sc_hd__o21ba_2
X_9206_ _9220_/CLK _9206_/D VGND VGND VPWR VPWR _9206_/Q sky130_fd_sc_hd__dfxtp_2
X_6418_ _6411_/X _6413_/Y _6414_/X _6417_/X VGND VGND VPWR VPWR _6464_/A sky130_fd_sc_hd__a211oi_1
X_9137_ _9214_/CLK _9137_/D VGND VGND VPWR VPWR _9137_/Q sky130_fd_sc_hd__dfxtp_1
X_7398_ _7539_/B _7539_/C _7539_/A VGND VGND VPWR VPWR _7398_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6349_ _6350_/A _6350_/B _6350_/C VGND VGND VPWR VPWR _6372_/B sky130_fd_sc_hd__a21oi_1
XFILLER_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9068_ _9090_/CLK _9068_/D VGND VGND VPWR VPWR _9068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8019_ _8128_/B _8019_/B VGND VGND VPWR VPWR _8025_/A sky130_fd_sc_hd__or2_1
XFILLER_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5720_ _5765_/A _4891_/X _4535_/X VGND VGND VPWR VPWR _5720_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5651_ _5583_/X _5650_/X _5674_/S VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8370_ _8370_/A _8370_/B VGND VGND VPWR VPWR _8373_/A sky130_fd_sc_hd__nor2_1
X_5582_ _5754_/B _5510_/X _5511_/X _5580_/X _5581_/X VGND VGND VPWR VPWR _9142_/D
+ sky130_fd_sc_hd__o221a_2
X_4602_ _5509_/A _4602_/B VGND VGND VPWR VPWR _4602_/Y sky130_fd_sc_hd__nor2_1
X_4533_ _9121_/Q _9113_/Q VGND VGND VPWR VPWR _4691_/A sky130_fd_sc_hd__xor2_4
X_7321_ _7321_/A _7321_/B VGND VGND VPWR VPWR _7321_/X sky130_fd_sc_hd__or2_1
X_7252_ _5908_/B _7119_/C _9183_/Q _6998_/A VGND VGND VPWR VPWR _7252_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6203_ _6204_/A _6204_/B _6204_/C VGND VGND VPWR VPWR _6292_/A sky130_fd_sc_hd__a21oi_2
X_7183_ _7406_/A _7552_/A _7182_/Y VGND VGND VPWR VPWR _7290_/A sky130_fd_sc_hd__a21bo_1
X_6134_ _6702_/B VGND VGND VPWR VPWR _7307_/B sky130_fd_sc_hd__clkbuf_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6065_ _9170_/Q VGND VGND VPWR VPWR _7148_/B sky130_fd_sc_hd__clkbuf_2
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5016_ _4641_/A _5015_/X _4961_/X VGND VGND VPWR VPWR _5017_/B sky130_fd_sc_hd__o21a_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6967_ _7531_/A _8844_/A _8733_/D _6875_/A VGND VGND VPWR VPWR _6986_/A sky130_fd_sc_hd__a22o_1
X_8706_ _8705_/A _8705_/B _8705_/C VGND VGND VPWR VPWR _8768_/A sky130_fd_sc_hd__a21oi_2
XFILLER_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5918_ _5918_/A _5918_/B _5918_/C VGND VGND VPWR VPWR _5930_/B sky130_fd_sc_hd__nand3_2
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6898_ _6791_/A _6790_/B _6790_/A VGND VGND VPWR VPWR _6993_/A sky130_fd_sc_hd__o21ba_1
X_8637_ _8637_/A _8637_/B VGND VGND VPWR VPWR _8639_/C sky130_fd_sc_hd__and2_1
X_5849_ _9165_/Q _6447_/A _6055_/A _6025_/A VGND VGND VPWR VPWR _5854_/A sky130_fd_sc_hd__and4_1
X_8568_ _8568_/A _8816_/B VGND VGND VPWR VPWR _8569_/B sky130_fd_sc_hd__nand2_1
X_7519_ _7658_/B _7517_/X _7518_/C _7518_/Y VGND VGND VPWR VPWR _7521_/A sky130_fd_sc_hd__o211a_1
X_8499_ _8499_/A _8499_/B VGND VGND VPWR VPWR _8501_/C sky130_fd_sc_hd__or2_1
XFILLER_103_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7870_ _8071_/A _8069_/A _8156_/C _8154_/B VGND VGND VPWR VPWR _7870_/X sky130_fd_sc_hd__and4_1
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6821_ _7822_/C VGND VGND VPWR VPWR _7938_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_63_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6752_ _6752_/A _6687_/B VGND VGND VPWR VPWR _6767_/B sky130_fd_sc_hd__or2b_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6683_ _8038_/A _7485_/A _6684_/C VGND VGND VPWR VPWR _6751_/B sky130_fd_sc_hd__a21oi_1
X_5703_ _5393_/A _4847_/X _4585_/A VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__a21o_1
X_8422_ _8422_/A _8422_/B VGND VGND VPWR VPWR _8423_/C sky130_fd_sc_hd__xor2_1
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5634_ _5634_/A _5634_/B VGND VGND VPWR VPWR _5634_/Y sky130_fd_sc_hd__nand2_1
X_8353_ _8245_/Y _8249_/B _8522_/A _8154_/X VGND VGND VPWR VPWR _8355_/B sky130_fd_sc_hd__a2bb2o_1
X_7304_ _7804_/A _8052_/B _7202_/A _7200_/B VGND VGND VPWR VPWR _7312_/A sky130_fd_sc_hd__a31o_1
X_5565_ _5003_/X _5119_/A _4597_/A VGND VGND VPWR VPWR _5565_/Y sky130_fd_sc_hd__a21oi_1
X_8284_ _8410_/B _8284_/B VGND VGND VPWR VPWR _8286_/A sky130_fd_sc_hd__xnor2_1
X_5496_ _5394_/X _5129_/X _5175_/X VGND VGND VPWR VPWR _5496_/Y sky130_fd_sc_hd__a21oi_1
X_7235_ _7235_/A _7235_/B _7235_/C VGND VGND VPWR VPWR _7235_/Y sky130_fd_sc_hd__nand3_2
X_7166_ _7166_/A _7166_/B _7218_/A VGND VGND VPWR VPWR _7274_/B sky130_fd_sc_hd__or3_2
XFILLER_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6117_ _6118_/B _6118_/C _6118_/A VGND VGND VPWR VPWR _6119_/A sky130_fd_sc_hd__a21oi_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7097_/A _7097_/B VGND VGND VPWR VPWR _7099_/B sky130_fd_sc_hd__xnor2_1
XFILLER_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6048_ _6048_/A VGND VGND VPWR VPWR _6125_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7999_ _7890_/A _7890_/B _7889_/B VGND VGND VPWR VPWR _8001_/B sky130_fd_sc_hd__o21a_1
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5350_ _5169_/A _5124_/A _4672_/A VGND VGND VPWR VPWR _5350_/Y sky130_fd_sc_hd__a21oi_1
X_5281_ _5120_/X _5280_/X _5281_/S VGND VGND VPWR VPWR _5281_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7020_ _7020_/A _7020_/B VGND VGND VPWR VPWR _7021_/B sky130_fd_sc_hd__nor2_1
XFILLER_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8971_ _8775_/B _8880_/Y _8967_/Y _8970_/Y VGND VGND VPWR VPWR _8972_/B sky130_fd_sc_hd__a31oi_4
X_7922_ _8177_/A _8269_/A _8175_/D _8038_/A VGND VGND VPWR VPWR _7924_/A sky130_fd_sc_hd__a22oi_1
XFILLER_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7853_ _7853_/A _7853_/B VGND VGND VPWR VPWR _7855_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7784_ _7784_/A _7784_/B _7784_/C VGND VGND VPWR VPWR _7786_/A sky130_fd_sc_hd__or3_1
X_6804_ _6805_/A _6805_/B _6805_/C VGND VGND VPWR VPWR _6934_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4996_ _5052_/B VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6735_ _6837_/A _6735_/B VGND VGND VPWR VPWR _6737_/C sky130_fd_sc_hd__nand2_1
X_6666_ _7118_/A _7116_/D VGND VGND VPWR VPWR _6671_/A sky130_fd_sc_hd__nand2_1
X_8405_ _8405_/A _8405_/B _8412_/B VGND VGND VPWR VPWR _8405_/X sky130_fd_sc_hd__or3_2
X_6597_ _6597_/A _6597_/B VGND VGND VPWR VPWR _6599_/A sky130_fd_sc_hd__xnor2_1
X_5617_ _5339_/A _5170_/X _5615_/X _5616_/Y _5173_/X VGND VGND VPWR VPWR _5617_/X
+ sky130_fd_sc_hd__a221o_1
X_8336_ _8336_/A _8336_/B VGND VGND VPWR VPWR _8336_/X sky130_fd_sc_hd__or2_1
X_5548_ _4573_/X _5126_/X _5181_/X VGND VGND VPWR VPWR _5548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8267_ _8267_/A _8267_/B VGND VGND VPWR VPWR _8405_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5479_ _5364_/X _5478_/X _5552_/S VGND VGND VPWR VPWR _5479_/X sky130_fd_sc_hd__mux2_1
X_7218_ _7218_/A VGND VGND VPWR VPWR _7274_/A sky130_fd_sc_hd__inv_2
X_8198_ _8197_/A _8197_/B _8196_/Y VGND VGND VPWR VPWR _8199_/B sky130_fd_sc_hd__o21bai_2
X_7149_ _7149_/A _7149_/B VGND VGND VPWR VPWR _7150_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4850_ _5286_/A _4850_/B VGND VGND VPWR VPWR _4850_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6520_ _7037_/A VGND VGND VPWR VPWR _7694_/A sky130_fd_sc_hd__clkbuf_2
X_4781_ _4935_/A _4773_/Y _4787_/B _4940_/A _4783_/A VGND VGND VPWR VPWR _4781_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6451_ _6451_/A _6451_/B VGND VGND VPWR VPWR _6452_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9170_ _9210_/CLK _9170_/D VGND VGND VPWR VPWR _9170_/Q sky130_fd_sc_hd__dfxtp_4
X_5402_ _5402_/A VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__clkbuf_2
X_6382_ _6480_/B _6382_/B VGND VGND VPWR VPWR _6383_/B sky130_fd_sc_hd__xnor2_2
X_8121_ _8132_/A _8132_/B VGND VGND VPWR VPWR _8125_/A sky130_fd_sc_hd__xnor2_1
X_5333_ _5117_/A _5331_/X _5575_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8052_ _8175_/B _8052_/B VGND VGND VPWR VPWR _8053_/B sky130_fd_sc_hd__nand2_1
X_5264_ _5165_/X _5555_/A _4607_/A VGND VGND VPWR VPWR _5264_/Y sky130_fd_sc_hd__a21oi_1
X_7003_ _7003_/A _7134_/B VGND VGND VPWR VPWR _7110_/A sky130_fd_sc_hd__nor2_1
X_5195_ _4739_/X _5194_/X _4980_/A VGND VGND VPWR VPWR _5195_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8954_ _8954_/A _8954_/B VGND VGND VPWR VPWR _8955_/B sky130_fd_sc_hd__nand2_1
X_7905_ _7903_/X _8018_/A VGND VGND VPWR VPWR _7911_/B sky130_fd_sc_hd__and2b_1
X_8885_ _8885_/A _8921_/B VGND VGND VPWR VPWR _8886_/A sky130_fd_sc_hd__and2_1
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7836_ _7837_/B _7837_/C _7837_/A VGND VGND VPWR VPWR _7841_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7767_ _7767_/A _8720_/B _7767_/C VGND VGND VPWR VPWR _7876_/A sky130_fd_sc_hd__and3_1
X_4979_ _4944_/A _5093_/A _4739_/A VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__o21a_1
X_7698_ _7804_/A _7810_/B _7569_/D _7567_/X VGND VGND VPWR VPWR _7699_/B sky130_fd_sc_hd__a31o_1
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6718_ _6716_/C _6716_/Y _6714_/Y _6715_/X VGND VGND VPWR VPWR _6740_/C sky130_fd_sc_hd__o211ai_4
X_6649_ _6649_/A _6649_/B _6649_/C VGND VGND VPWR VPWR _6651_/A sky130_fd_sc_hd__or3_1
X_8319_ _8318_/A _8318_/B _8317_/Y VGND VGND VPWR VPWR _8423_/A sky130_fd_sc_hd__o21ba_1
XFILLER_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5951_ _5951_/A _5951_/B VGND VGND VPWR VPWR _5952_/B sky130_fd_sc_hd__and2_1
XFILLER_18_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8670_ _8670_/A _8670_/B VGND VGND VPWR VPWR _8671_/B sky130_fd_sc_hd__nor2_1
X_4902_ _9125_/Q _9117_/Q VGND VGND VPWR VPWR _4991_/A sky130_fd_sc_hd__nand2_1
X_5882_ _5886_/A _5886_/B VGND VGND VPWR VPWR _5885_/C sky130_fd_sc_hd__or2_1
XFILLER_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7621_ _7621_/A _7621_/B _7621_/C VGND VGND VPWR VPWR _7622_/B sky130_fd_sc_hd__nand3_4
X_4833_ _4833_/A _4937_/A VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__or2_2
X_7552_ _7552_/A _7552_/B VGND VGND VPWR VPWR _7552_/Y sky130_fd_sc_hd__nand2_1
X_4764_ _4929_/A _4924_/A VGND VGND VPWR VPWR _4764_/X sky130_fd_sc_hd__or2_2
X_7483_ _7610_/D VGND VGND VPWR VPWR _7959_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6503_ _7187_/A _7608_/A VGND VGND VPWR VPWR _6504_/B sky130_fd_sc_hd__nand2_1
X_9222_ _9222_/CLK _9222_/D VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
X_6434_ _6434_/A _6434_/B VGND VGND VPWR VPWR _6458_/B sky130_fd_sc_hd__nand2_1
X_4695_ _4739_/A VGND VGND VPWR VPWR _4891_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9153_ _9214_/CLK _9153_/D VGND VGND VPWR VPWR _9153_/Q sky130_fd_sc_hd__dfxtp_1
X_6365_ _6414_/B _6365_/B VGND VGND VPWR VPWR _6417_/C sky130_fd_sc_hd__xnor2_1
X_8104_ _8102_/X _7975_/B _8100_/Y _8203_/A VGND VGND VPWR VPWR _8203_/B sky130_fd_sc_hd__o211ai_4
XFILLER_88_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6296_ _6380_/A _6380_/B VGND VGND VPWR VPWR _6385_/B sky130_fd_sc_hd__xnor2_2
X_5316_ _5316_/A _5369_/A VGND VGND VPWR VPWR _5316_/Y sky130_fd_sc_hd__nand2_1
X_9084_ _9090_/CLK _9084_/D VGND VGND VPWR VPWR _9084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8035_ _8279_/A _8595_/C _8595_/D _8177_/A VGND VGND VPWR VPWR _8037_/A sky130_fd_sc_hd__a22oi_1
X_5247_ _5410_/A VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold15 hold2/X VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5178_ _9081_/Q VGND VGND VPWR VPWR _5179_/A sky130_fd_sc_hd__clkinv_2
XFILLER_56_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8937_ _8937_/A _8937_/B _8937_/C VGND VGND VPWR VPWR _8985_/A sky130_fd_sc_hd__nor3_1
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8868_ _8868_/A _8868_/B VGND VGND VPWR VPWR _8870_/B sky130_fd_sc_hd__xor2_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8799_ _8800_/A _8800_/B VGND VGND VPWR VPWR _8801_/A sky130_fd_sc_hd__or2_1
X_7819_ _8038_/A _8052_/B _7819_/C VGND VGND VPWR VPWR _7828_/B sky130_fd_sc_hd__and3_1
XFILLER_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6150_ _7327_/B VGND VGND VPWR VPWR _7706_/B sky130_fd_sc_hd__buf_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5043_/A _5100_/Y _5785_/S VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__mux2_2
X_6081_ _6081_/A _6081_/B VGND VGND VPWR VPWR _6085_/A sky130_fd_sc_hd__nor2_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/A _5032_/B VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__xnor2_1
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6983_ _6864_/A _6864_/B _6982_/X VGND VGND VPWR VPWR _6984_/B sky130_fd_sc_hd__a21bo_1
X_8722_ _8722_/A _8787_/A VGND VGND VPWR VPWR _8724_/C sky130_fd_sc_hd__nor2_1
X_5934_ _5952_/A _5951_/A _6000_/A _5932_/X VGND VGND VPWR VPWR _6047_/A sky130_fd_sc_hd__or4bb_4
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8653_ _8652_/B _8772_/A _8773_/A VGND VGND VPWR VPWR _8714_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5865_ _5898_/C _5865_/B VGND VGND VPWR VPWR _5952_/A sky130_fd_sc_hd__xnor2_2
X_7604_ _7730_/A _7604_/B _7604_/C _7604_/D VGND VGND VPWR VPWR _7605_/B sky130_fd_sc_hd__and4_1
X_4816_ _4816_/A _4816_/B VGND VGND VPWR VPWR _4828_/C sky130_fd_sc_hd__xor2_2
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8584_ _8584_/A VGND VGND VPWR VPWR _8716_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5796_ _6778_/B VGND VGND VPWR VPWR _7766_/A sky130_fd_sc_hd__clkbuf_4
X_7535_ _7535_/A _7535_/B VGND VGND VPWR VPWR _7536_/B sky130_fd_sc_hd__nor2_1
X_4747_ _4747_/A VGND VGND VPWR VPWR _9153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7466_ _7610_/C VGND VGND VPWR VPWR _8190_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4678_ _4982_/A _4897_/A VGND VGND VPWR VPWR _5511_/A sky130_fd_sc_hd__nand2_2
X_9205_ _9214_/CLK _9205_/D VGND VGND VPWR VPWR _9205_/Q sky130_fd_sc_hd__dfxtp_2
X_6417_ _6875_/A _8438_/A _6417_/C VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and3_1
X_7397_ _7397_/A _7397_/B VGND VGND VPWR VPWR _7539_/A sky130_fd_sc_hd__xnor2_1
X_9136_ _9222_/CLK _9136_/D VGND VGND VPWR VPWR _9136_/Q sky130_fd_sc_hd__dfxtp_1
X_6348_ _6248_/A _6332_/B _6248_/C _6263_/X VGND VGND VPWR VPWR _6350_/C sky130_fd_sc_hd__a31o_1
XFILLER_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6279_ _6279_/A _6279_/B VGND VGND VPWR VPWR _6280_/B sky130_fd_sc_hd__nor2_1
X_9067_ _9199_/CLK _9067_/D VGND VGND VPWR VPWR _9067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8018_ _8018_/A _8018_/B _8018_/C VGND VGND VPWR VPWR _8019_/B sky130_fd_sc_hd__and3_1
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_5650_ _5633_/Y _5649_/Y _5281_/S _5754_/B VGND VGND VPWR VPWR _5650_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4601_ _4870_/S _4594_/X _4636_/A VGND VGND VPWR VPWR _4602_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5581_ _5581_/A _5604_/B VGND VGND VPWR VPWR _5581_/X sky130_fd_sc_hd__or2_1
X_7320_ _7319_/A _7319_/B _7319_/C VGND VGND VPWR VPWR _7533_/A sky130_fd_sc_hd__a21oi_2
XFILLER_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7251_ _7251_/A _7251_/B VGND VGND VPWR VPWR _7265_/B sky130_fd_sc_hd__nand2_1
X_6202_ _6202_/A _6282_/A VGND VGND VPWR VPWR _6204_/C sky130_fd_sc_hd__or2_1
X_7182_ _7182_/A _7182_/B VGND VGND VPWR VPWR _7182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6133_ _7006_/A VGND VGND VPWR VPWR _7770_/A sky130_fd_sc_hd__clkbuf_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6064_ _6223_/A _6572_/B _6925_/A _6325_/B VGND VGND VPWR VPWR _6068_/C sky130_fd_sc_hd__a22o_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5015_ _5132_/A _5014_/X _4958_/X VGND VGND VPWR VPWR _5015_/X sky130_fd_sc_hd__o21a_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6966_ _8595_/D VGND VGND VPWR VPWR _8733_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_81_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8705_ _8705_/A _8705_/B _8705_/C VGND VGND VPWR VPWR _8705_/X sky130_fd_sc_hd__and3_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5917_ _5918_/A _5918_/B _5918_/C VGND VGND VPWR VPWR _5930_/A sky130_fd_sc_hd__a21o_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6897_ _6897_/A _6897_/B VGND VGND VPWR VPWR _6899_/A sky130_fd_sc_hd__xnor2_1
X_8636_ _8635_/A _8635_/B _8634_/Y VGND VGND VPWR VPWR _8637_/B sky130_fd_sc_hd__o21bai_2
X_5848_ _9196_/Q VGND VGND VPWR VPWR _6447_/A sky130_fd_sc_hd__clkbuf_2
X_8567_ _8567_/A _8567_/B VGND VGND VPWR VPWR _8569_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5779_ _4636_/A _5778_/Y _4876_/A VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__o21a_1
X_7518_ _7518_/A _7518_/B _7518_/C VGND VGND VPWR VPWR _7518_/Y sky130_fd_sc_hd__nand3_2
X_8498_ _8498_/A _8909_/B _8498_/C VGND VGND VPWR VPWR _8499_/B sky130_fd_sc_hd__and3_1
X_7449_ _7449_/A _7449_/B VGND VGND VPWR VPWR _7449_/X sky130_fd_sc_hd__or2_1
XFILLER_103_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9119_ _9221_/CLK _9191_/Q VGND VGND VPWR VPWR _9119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6820_ _9208_/Q VGND VGND VPWR VPWR _7822_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6751_ _6751_/A _6751_/B _6805_/B VGND VGND VPWR VPWR _6767_/A sky130_fd_sc_hd__or3_2
XFILLER_50_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6682_ _6805_/A _6682_/B VGND VGND VPWR VPWR _6684_/C sky130_fd_sc_hd__nor2_1
X_5702_ _5389_/A _5369_/A _5701_/X VGND VGND VPWR VPWR _5702_/Y sky130_fd_sc_hd__a21oi_1
X_8421_ _8421_/A _8325_/X VGND VGND VPWR VPWR _8422_/B sky130_fd_sc_hd__or2b_1
X_5633_ _5534_/A _4889_/A _4737_/X VGND VGND VPWR VPWR _5633_/Y sky130_fd_sc_hd__a21oi_1
X_8352_ _8352_/A _8352_/B VGND VGND VPWR VPWR _8355_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5564_ _5215_/X _5194_/A _5562_/X _5563_/Y _5058_/A VGND VGND VPWR VPWR _5564_/X
+ sky130_fd_sc_hd__a221o_1
X_7303_ _7569_/C VGND VGND VPWR VPWR _7804_/A sky130_fd_sc_hd__clkbuf_2
X_8283_ _8176_/A _8179_/B _8176_/B VGND VGND VPWR VPWR _8284_/B sky130_fd_sc_hd__o21ba_1
X_5495_ _5266_/X _5116_/A _5493_/X _5494_/Y _5173_/X VGND VGND VPWR VPWR _5495_/X
+ sky130_fd_sc_hd__a221o_1
X_7234_ _7234_/A _7234_/B VGND VGND VPWR VPWR _7235_/C sky130_fd_sc_hd__nand2_1
X_7165_ _7166_/B _7218_/A _7166_/A VGND VGND VPWR VPWR _7165_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6294_/A _6116_/B VGND VGND VPWR VPWR _6118_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/A _7696_/B VGND VGND VPWR VPWR _7097_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6047_ _6047_/A _6047_/B _6131_/A _6047_/D VGND VGND VPWR VPWR _6048_/A sky130_fd_sc_hd__or4_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7998_ _8081_/A _7998_/B VGND VGND VPWR VPWR _8001_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6949_ _6949_/A _6949_/B VGND VGND VPWR VPWR _6959_/B sky130_fd_sc_hd__xnor2_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8619_ _8619_/A _8619_/B VGND VGND VPWR VPWR _8620_/B sky130_fd_sc_hd__or2_1
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5280_ _5187_/X _5206_/X _5275_/X _5279_/Y VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8970_ _8970_/A VGND VGND VPWR VPWR _8970_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7921_ _7923_/B VGND VGND VPWR VPWR _8177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7852_ _7852_/A _8243_/A _7852_/C _8148_/A VGND VGND VPWR VPWR _7853_/B sky130_fd_sc_hd__and4_1
XFILLER_51_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7783_ _7783_/A _7783_/B VGND VGND VPWR VPWR _7784_/C sky130_fd_sc_hd__xor2_1
X_6803_ _6919_/A _6803_/B VGND VGND VPWR VPWR _6805_/C sky130_fd_sc_hd__xnor2_1
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4995_ _4995_/A _5033_/B VGND VGND VPWR VPWR _5052_/B sky130_fd_sc_hd__nor2_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6734_ _6734_/A _6734_/B VGND VGND VPWR VPWR _6735_/B sky130_fd_sc_hd__or2_1
X_8404_ _8403_/B _8494_/B _8403_/A VGND VGND VPWR VPWR _8404_/Y sky130_fd_sc_hd__a21oi_2
X_6665_ _6665_/A _6665_/B VGND VGND VPWR VPWR _6774_/A sky130_fd_sc_hd__xnor2_1
X_6596_ _6596_/A _6596_/B VGND VGND VPWR VPWR _6597_/B sky130_fd_sc_hd__nor2_1
X_5616_ _5558_/X _5132_/X _5414_/X VGND VGND VPWR VPWR _5616_/Y sky130_fd_sc_hd__a21oi_1
X_8335_ _8335_/A _8335_/B VGND VGND VPWR VPWR _9097_/D sky130_fd_sc_hd__xor2_1
X_5547_ _5315_/A _5177_/X _5545_/X _5546_/Y _5126_/A VGND VGND VPWR VPWR _5547_/X
+ sky130_fd_sc_hd__a221o_1
X_8266_ _8266_/A _8266_/B VGND VGND VPWR VPWR _8267_/B sky130_fd_sc_hd__nand2_2
X_5478_ _5339_/X _5477_/X _5575_/S VGND VGND VPWR VPWR _5478_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7217_ _7215_/Y _7103_/B _7213_/X _7394_/A VGND VGND VPWR VPWR _7394_/B sky130_fd_sc_hd__a211oi_4
X_8197_ _8197_/A _8197_/B _8196_/Y VGND VGND VPWR VPWR _8199_/A sky130_fd_sc_hd__or3b_1
XFILLER_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_7148_ _7148_/A _7148_/B _7222_/C _7148_/D VGND VGND VPWR VPWR _7149_/B sky130_fd_sc_hd__and4_1
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7079_ _7079_/A _7079_/B VGND VGND VPWR VPWR _7087_/A sky130_fd_sc_hd__or2_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4780_ _4780_/A VGND VGND VPWR VPWR _4940_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6450_ _7506_/A _7042_/C _7822_/B _5818_/X VGND VGND VPWR VPWR _6451_/B sky130_fd_sc_hd__a22oi_1
X_5401_ _5364_/X _5365_/X _5366_/X _5399_/X _5400_/X VGND VGND VPWR VPWR _9135_/D
+ sky130_fd_sc_hd__o221a_4
X_6381_ _6385_/A _6385_/B _6480_/A VGND VGND VPWR VPWR _6382_/B sky130_fd_sc_hd__o21a_1
X_8120_ _8131_/A _8120_/B VGND VGND VPWR VPWR _8132_/B sky130_fd_sc_hd__xnor2_1
X_5332_ _5739_/S VGND VGND VPWR VPWR _5575_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8051_ _8051_/A _8051_/B VGND VGND VPWR VPWR _8053_/A sky130_fd_sc_hd__nor2_1
X_5263_ _9079_/Q VGND VGND VPWR VPWR _5555_/A sky130_fd_sc_hd__clkbuf_4
X_7002_ _7134_/A _7000_/Y _7361_/C _7610_/C VGND VGND VPWR VPWR _7134_/B sky130_fd_sc_hd__and4bb_1
X_5194_ _5194_/A VGND VGND VPWR VPWR _5194_/X sky130_fd_sc_hd__buf_4
XFILLER_83_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8953_ _8954_/A _8954_/B VGND VGND VPWR VPWR _8955_/A sky130_fd_sc_hd__or2_1
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7904_ _7903_/A _7903_/B _7903_/C VGND VGND VPWR VPWR _8018_/A sky130_fd_sc_hd__a21o_1
X_8884_ _8966_/A _8884_/B VGND VGND VPWR VPWR _8921_/B sky130_fd_sc_hd__nand2_1
X_7835_ _7745_/A _7745_/B _7745_/C VGND VGND VPWR VPWR _7837_/A sky130_fd_sc_hd__a21bo_1
XFILLER_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7766_ _7766_/A _8720_/B VGND VGND VPWR VPWR _7984_/A sky130_fd_sc_hd__nand2_1
X_4978_ _5696_/S _4974_/X _4976_/X _4977_/X VGND VGND VPWR VPWR _4978_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7697_ _7697_/A _7697_/B VGND VGND VPWR VPWR _7699_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6717_ _6714_/Y _6715_/X _6716_/C _6716_/Y VGND VGND VPWR VPWR _6740_/B sky130_fd_sc_hd__a211o_1
XFILLER_50_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6648_ _6655_/C _6648_/B VGND VGND VPWR VPWR _6649_/C sky130_fd_sc_hd__xor2_1
X_8318_ _8318_/A _8318_/B _8317_/Y VGND VGND VPWR VPWR _8320_/A sky130_fd_sc_hd__nor3b_1
X_6579_ _6579_/A _6579_/B VGND VGND VPWR VPWR _6580_/C sky130_fd_sc_hd__xnor2_1
XFILLER_105_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8249_ _8249_/A _8249_/B VGND VGND VPWR VPWR _8251_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5950_ _9056_/A _9060_/B VGND VGND VPWR VPWR _9057_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4901_ _4901_/A VGND VGND VPWR VPWR _4905_/A sky130_fd_sc_hd__clkinv_2
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7620_ _7621_/B _7621_/C _7621_/A VGND VGND VPWR VPWR _7622_/A sky130_fd_sc_hd__a21o_1
X_5881_ _5881_/A _5892_/A VGND VGND VPWR VPWR _5886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4832_ _4837_/A _4943_/A VGND VGND VPWR VPWR _4937_/A sky130_fd_sc_hd__nor2_1
X_7551_ _7408_/A _7408_/C _7549_/A _7550_/X _7553_/B VGND VGND VPWR VPWR _7677_/B
+ sky130_fd_sc_hd__a311oi_4
X_4763_ _4837_/A _4960_/A VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__nor2_1
X_7482_ _7482_/A _7482_/B VGND VGND VPWR VPWR _7600_/A sky130_fd_sc_hd__nor2_1
X_4694_ _9110_/Q VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__clkbuf_2
X_6502_ _6502_/A _6502_/B VGND VGND VPWR VPWR _6504_/A sky130_fd_sc_hd__nor2_1
X_9221_ _9221_/CLK _9221_/D VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
X_6433_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6458_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9152_ _9213_/CLK _9152_/D VGND VGND VPWR VPWR _9152_/Q sky130_fd_sc_hd__dfxtp_1
X_6364_ _6280_/A _6279_/B _6279_/A VGND VGND VPWR VPWR _6365_/B sky130_fd_sc_hd__o21ba_1
X_8103_ _8100_/Y _8203_/A _8102_/X _7975_/B VGND VGND VPWR VPWR _8105_/B sky130_fd_sc_hd__a211o_1
XFILLER_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5315_ _5315_/A VGND VGND VPWR VPWR _5315_/X sky130_fd_sc_hd__clkbuf_2
X_6295_ _6294_/Y _6211_/A _6211_/B VGND VGND VPWR VPWR _6380_/B sky130_fd_sc_hd__o21ba_1
X_9083_ _9090_/CLK _9083_/D VGND VGND VPWR VPWR _9083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8034_ _8036_/B VGND VGND VPWR VPWR _8279_/A sky130_fd_sc_hd__clkbuf_2
X_5246_ _9080_/Q VGND VGND VPWR VPWR _5246_/Y sky130_fd_sc_hd__inv_2
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__buf_2
X_5177_ _5177_/A VGND VGND VPWR VPWR _5177_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8936_ _8936_/A _8936_/B VGND VGND VPWR VPWR _8937_/C sky130_fd_sc_hd__or2_1
X_8867_ _8867_/A _8867_/B VGND VGND VPWR VPWR _8868_/B sky130_fd_sc_hd__nand2_1
X_8798_ _8867_/A _8798_/B VGND VGND VPWR VPWR _8800_/B sky130_fd_sc_hd__and2_1
X_7818_ _7710_/A _7818_/B VGND VGND VPWR VPWR _7830_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7749_ _8150_/C VGND VGND VPWR VPWR _8464_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6080_ _6500_/B _6151_/A _6778_/B _7453_/A VGND VGND VPWR VPWR _6081_/B sky130_fd_sc_hd__and4_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5100_ _5676_/B _5043_/Y _5099_/X VGND VGND VPWR VPWR _5100_/Y sky130_fd_sc_hd__a21oi_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B VGND VGND VPWR VPWR _5032_/B sky130_fd_sc_hd__nor2_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8721_ _8721_/A _8721_/B _8887_/A VGND VGND VPWR VPWR _8787_/A sky130_fd_sc_hd__and3_1
XFILLER_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6982_ _6982_/A _6863_/B VGND VGND VPWR VPWR _6982_/X sky130_fd_sc_hd__or2b_1
XFILLER_80_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5933_ _5952_/A _5951_/A _6000_/A _5932_/X VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8652_ _8773_/A _8652_/B _8772_/A VGND VGND VPWR VPWR _8652_/X sky130_fd_sc_hd__and3_1
X_5864_ _5862_/X _5898_/B VGND VGND VPWR VPWR _5865_/B sky130_fd_sc_hd__and2b_1
X_8583_ _8522_/A _8523_/A _8522_/B VGND VGND VPWR VPWR _8592_/B sky130_fd_sc_hd__o21bai_2
X_7603_ _8050_/A _7847_/A _7459_/D _7730_/A VGND VGND VPWR VPWR _7605_/A sky130_fd_sc_hd__a22oi_1
X_4815_ _4901_/A _4815_/B VGND VGND VPWR VPWR _4816_/B sky130_fd_sc_hd__nand2_2
X_5795_ _5908_/B VGND VGND VPWR VPWR _6778_/B sky130_fd_sc_hd__buf_2
X_7534_ _7533_/A _7533_/B _7532_/Y VGND VGND VPWR VPWR _7535_/B sky130_fd_sc_hd__o21ba_1
X_4746_ _4966_/B _4744_/Y _5653_/B VGND VGND VPWR VPWR _4747_/A sky130_fd_sc_hd__mux2_4
X_7465_ _7465_/A VGND VGND VPWR VPWR _8050_/B sky130_fd_sc_hd__clkbuf_2
X_4677_ _4677_/A _4677_/B _4677_/C VGND VGND VPWR VPWR _4897_/A sky130_fd_sc_hd__or3_2
X_9204_ _9210_/CLK _9204_/D VGND VGND VPWR VPWR _9204_/Q sky130_fd_sc_hd__dfxtp_2
X_6416_ _8587_/A VGND VGND VPWR VPWR _8438_/A sky130_fd_sc_hd__buf_4
X_7396_ _7396_/A _7396_/B VGND VGND VPWR VPWR _7397_/B sky130_fd_sc_hd__nor2_1
X_9135_ _9222_/CLK _9135_/D VGND VGND VPWR VPWR _9135_/Q sky130_fd_sc_hd__dfxtp_1
X_6347_ _6347_/A _6347_/B _6347_/C VGND VGND VPWR VPWR _6350_/B sky130_fd_sc_hd__nand3_1
XFILLER_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9066_ _9224_/CLK hold9/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
X_6278_ _6700_/A _7852_/A _8243_/A _6359_/A VGND VGND VPWR VPWR _6279_/B sky130_fd_sc_hd__a22oi_2
XFILLER_69_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8017_ _8018_/A _8018_/B _8018_/C VGND VGND VPWR VPWR _8128_/B sky130_fd_sc_hd__a21oi_1
X_5229_ _5169_/A _5581_/A _4548_/A VGND VGND VPWR VPWR _5229_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8919_ _8876_/A _8876_/B _8874_/B VGND VGND VPWR VPWR _8920_/B sky130_fd_sc_hd__a21o_1
XFILLER_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4600_ _4600_/A VGND VGND VPWR VPWR _4636_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5580_ _5534_/X _5579_/X _5603_/S VGND VGND VPWR VPWR _5580_/X sky130_fd_sc_hd__mux2_1
X_7250_ _7250_/A _7124_/A VGND VGND VPWR VPWR _7265_/A sky130_fd_sc_hd__or2b_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6201_ _6968_/A _6968_/B _8156_/A _8156_/B VGND VGND VPWR VPWR _6282_/A sky130_fd_sc_hd__and4_1
X_7181_ _7406_/A _7552_/A VGND VGND VPWR VPWR _9087_/D sky130_fd_sc_hd__xor2_1
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6132_ _6132_/A _6221_/B VGND VGND VPWR VPWR _6301_/A sky130_fd_sc_hd__nor2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6063_ _7259_/B VGND VGND VPWR VPWR _6325_/B sky130_fd_sc_hd__clkbuf_2
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5164_/A _5013_/X _4954_/Y VGND VGND VPWR VPWR _5014_/X sky130_fd_sc_hd__o21a_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6965_ _8175_/D VGND VGND VPWR VPWR _8595_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_81_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8704_ _8704_/A _8761_/B VGND VGND VPWR VPWR _8705_/C sky130_fd_sc_hd__or2_1
X_5916_ _5861_/A _5860_/B _5858_/X VGND VGND VPWR VPWR _5918_/C sky130_fd_sc_hd__a21o_1
X_6896_ _6896_/A _6896_/B VGND VGND VPWR VPWR _6897_/B sky130_fd_sc_hd__nor2_1
X_8635_ _8635_/A _8635_/B _8634_/Y VGND VGND VPWR VPWR _8637_/A sky130_fd_sc_hd__or3b_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5847_ _5847_/A _5847_/B VGND VGND VPWR VPWR _5861_/A sky130_fd_sc_hd__xnor2_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8566_ _8565_/A _8565_/B _8564_/Y VGND VGND VPWR VPWR _8567_/B sky130_fd_sc_hd__o21ba_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5778_ _5621_/X _5777_/Y _4874_/S VGND VGND VPWR VPWR _5778_/Y sky130_fd_sc_hd__a21oi_1
X_7517_ _7516_/B _7658_/A _7516_/A VGND VGND VPWR VPWR _7517_/X sky130_fd_sc_hd__o21a_1
X_8497_ _8498_/A _8756_/B _8498_/C VGND VGND VPWR VPWR _8499_/A sky130_fd_sc_hd__a21oi_1
X_4729_ _5736_/S VGND VGND VPWR VPWR _5692_/S sky130_fd_sc_hd__clkbuf_2
X_7448_ _7447_/A _7447_/B _7447_/C VGND VGND VPWR VPWR _7559_/A sky130_fd_sc_hd__a21oi_2
X_7379_ _7377_/C _7377_/Y _7375_/X _7376_/Y VGND VGND VPWR VPWR _7379_/X sky130_fd_sc_hd__a211o_2
XFILLER_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9118_ _9218_/CLK hold1/X VGND VGND VPWR VPWR _9118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9049_ _9049_/A _9049_/B VGND VGND VPWR VPWR _9111_/D sky130_fd_sc_hd__xor2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6750_ _6750_/A _6745_/B VGND VGND VPWR VPWR _6848_/A sky130_fd_sc_hd__or2b_1
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5701_ _5313_/A _5420_/A _5146_/X _5194_/A _4856_/A VGND VGND VPWR VPWR _5701_/X
+ sky130_fd_sc_hd__a221o_1
X_6681_ _6424_/D _6143_/B _7706_/B _6907_/A VGND VGND VPWR VPWR _6682_/B sky130_fd_sc_hd__a22oi_1
X_8420_ _8420_/A _8420_/B VGND VGND VPWR VPWR _8422_/A sky130_fd_sc_hd__nor2_1
X_5632_ _5632_/A VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8351_ _8349_/X _8351_/B _8351_/C _8351_/D VGND VGND VPWR VPWR _8352_/B sky130_fd_sc_hd__and4b_1
X_5563_ _4862_/A _9086_/Q _5215_/A VGND VGND VPWR VPWR _5563_/Y sky130_fd_sc_hd__a21oi_1
X_7302_ _7302_/A _7302_/B VGND VGND VPWR VPWR _7449_/A sky130_fd_sc_hd__or2_1
X_8282_ _8282_/A _8282_/B VGND VGND VPWR VPWR _8410_/B sky130_fd_sc_hd__xnor2_1
X_5494_ _5382_/X _5389_/X _5414_/X VGND VGND VPWR VPWR _5494_/Y sky130_fd_sc_hd__a21oi_1
X_7233_ _7233_/A _7233_/B VGND VGND VPWR VPWR _7234_/B sky130_fd_sc_hd__nand2_1
X_7164_ _7164_/A _7164_/B VGND VGND VPWR VPWR _7166_/A sky130_fd_sc_hd__xnor2_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6875_/A _8349_/A _6107_/X _6108_/X VGND VGND VPWR VPWR _6116_/B sky130_fd_sc_hd__a211oi_1
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7095_ _9213_/Q VGND VGND VPWR VPWR _7696_/B sky130_fd_sc_hd__clkbuf_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6046_ _6047_/A _6047_/B _6131_/A _6047_/D VGND VGND VPWR VPWR _6049_/C sky130_fd_sc_hd__o22ai_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7997_ _7997_/A _7997_/B VGND VGND VPWR VPWR _7998_/B sky130_fd_sc_hd__nand2_1
X_6948_ _6948_/A _6948_/B VGND VGND VPWR VPWR _6949_/B sky130_fd_sc_hd__nor2_2
X_6879_ _6879_/A _6940_/B _6879_/C VGND VGND VPWR VPWR _6882_/C sky130_fd_sc_hd__nor3_1
X_8618_ _8619_/A _8619_/B VGND VGND VPWR VPWR _8620_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8549_ _8473_/A _8473_/B _8472_/B VGND VGND VPWR VPWR _8551_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7920_ _7920_/A _7920_/B VGND VGND VPWR VPWR _7952_/B sky130_fd_sc_hd__or2_1
XFILLER_48_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7851_ _8091_/B _7748_/A _8148_/A _8091_/A VGND VGND VPWR VPWR _7853_/A sky130_fd_sc_hd__a22oi_1
X_6802_ _6802_/A _6802_/B VGND VGND VPWR VPWR _6803_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7782_ _7782_/A _7899_/B VGND VGND VPWR VPWR _7783_/B sky130_fd_sc_hd__xnor2_4
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4994_ _4993_/B _4994_/B VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__and2b_1
X_6733_ _6734_/A _6734_/B VGND VGND VPWR VPWR _6837_/A sky130_fd_sc_hd__nand2_2
X_6664_ _6664_/A _6664_/B VGND VGND VPWR VPWR _6665_/B sky130_fd_sc_hd__nor2_1
X_8403_ _8403_/A _8403_/B _8494_/B VGND VGND VPWR VPWR _8490_/B sky130_fd_sc_hd__and3_2
X_5615_ _5287_/A _5165_/X _5613_/X _5614_/Y _4607_/A VGND VGND VPWR VPWR _5615_/X
+ sky130_fd_sc_hd__a221o_1
X_6595_ _6325_/A _6663_/C _7465_/A _5818_/X VGND VGND VPWR VPWR _6596_/B sky130_fd_sc_hd__a22oi_1
X_8334_ _8231_/A _8231_/B _8230_/A _8333_/Y VGND VGND VPWR VPWR _8335_/B sky130_fd_sc_hd__o31a_1
X_5546_ _5450_/X _5129_/X _5175_/X VGND VGND VPWR VPWR _5546_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8265_ _8266_/A _8266_/B VGND VGND VPWR VPWR _8267_/A sky130_fd_sc_hd__or2_1
X_5477_ _5315_/A _5476_/X _5527_/S VGND VGND VPWR VPWR _5477_/X sky130_fd_sc_hd__mux2_1
X_7216_ _7213_/X _7394_/A _7215_/Y _7103_/B VGND VGND VPWR VPWR _7277_/A sky130_fd_sc_hd__o211a_1
X_8196_ _8196_/A _8196_/B VGND VGND VPWR VPWR _8196_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ _7325_/A _7728_/B _7728_/D _6607_/A VGND VGND VPWR VPWR _7149_/A sky130_fd_sc_hd__a22oi_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _7078_/A _7078_/B VGND VGND VPWR VPWR _7088_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6029_ _6029_/A _6029_/B VGND VGND VPWR VPWR _6032_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5400_ _9073_/Q _5482_/B VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__or2_1
X_6380_ _6380_/A _6380_/B VGND VGND VPWR VPWR _6480_/A sky130_fd_sc_hd__or2_1
X_5331_ _5120_/A _5330_/X _5527_/S VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__mux2_1
X_8050_ _8050_/A _8050_/B _8050_/C _8050_/D VGND VGND VPWR VPWR _8051_/B sky130_fd_sc_hd__and4_1
X_7001_ _7767_/A _7847_/D _7134_/A _7000_/Y VGND VGND VPWR VPWR _7003_/A sky130_fd_sc_hd__o2bb2a_1
X_5262_ _5247_/X _5248_/Y _5259_/X _5261_/Y _4558_/A VGND VGND VPWR VPWR _5262_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5193_ _5205_/A VGND VGND VPWR VPWR _5194_/A sky130_fd_sc_hd__inv_2
XFILLER_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8952_ _8952_/A _8952_/B VGND VGND VPWR VPWR _8954_/B sky130_fd_sc_hd__nand2_1
X_7903_ _7903_/A _7903_/B _7903_/C VGND VGND VPWR VPWR _7903_/X sky130_fd_sc_hd__and3_1
X_8883_ _8966_/A _8884_/B VGND VGND VPWR VPWR _8885_/A sky130_fd_sc_hd__or2_1
X_7834_ _7834_/A _7834_/B VGND VGND VPWR VPWR _7837_/C sky130_fd_sc_hd__or2_1
XFILLER_24_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7765_ _8243_/B VGND VGND VPWR VPWR _8720_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4977_ _4737_/A _4940_/B _4940_/C _4739_/A VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__a31o_1
X_6716_ _6716_/A _6716_/B _6716_/C VGND VGND VPWR VPWR _6716_/Y sky130_fd_sc_hd__nor3_2
X_7696_ _7694_/X _7696_/B _7696_/C _7696_/D VGND VGND VPWR VPWR _7697_/B sky130_fd_sc_hd__and4b_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6647_ _6655_/A _6655_/B _6653_/A VGND VGND VPWR VPWR _6648_/B sky130_fd_sc_hd__a21o_1
X_6578_ _6693_/B _6578_/B VGND VGND VPWR VPWR _6579_/B sky130_fd_sc_hd__xnor2_1
X_8317_ _8322_/A _8933_/B _8183_/A _8316_/X VGND VGND VPWR VPWR _8317_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5529_ _5433_/X _5528_/X _5552_/S VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8248_ _8351_/C _8664_/C VGND VGND VPWR VPWR _8249_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8179_ _8179_/A _8179_/B VGND VGND VPWR VPWR _8316_/B sky130_fd_sc_hd__xnor2_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4900_ _4812_/X _4960_/B _4895_/X _4899_/Y VGND VGND VPWR VPWR _9155_/D sky130_fd_sc_hd__a2bb2o_4
X_5880_ _7689_/A _5945_/A VGND VGND VPWR VPWR _5886_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4831_ _4924_/A _4845_/B VGND VGND VPWR VPWR _4833_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4762_ _4762_/A VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__buf_2
X_7550_ _7553_/A _7550_/B VGND VGND VPWR VPWR _7550_/X sky130_fd_sc_hd__and2b_1
X_7481_ _7873_/A _8290_/A _7351_/B _7349_/X VGND VGND VPWR VPWR _7601_/A sky130_fd_sc_hd__a31o_1
X_6501_ _7419_/B _6927_/C _6361_/D _7201_/A VGND VGND VPWR VPWR _6502_/B sky130_fd_sc_hd__a22oi_2
X_4693_ _4837_/A _4842_/A VGND VGND VPWR VPWR _4693_/Y sky130_fd_sc_hd__nand2_4
X_9220_ _9220_/CLK _9220_/D VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_1
X_6432_ _6489_/A _6432_/B VGND VGND VPWR VPWR _6512_/A sky130_fd_sc_hd__xnor2_1
X_9151_ _9210_/CLK _9151_/D VGND VGND VPWR VPWR _9151_/Q sky130_fd_sc_hd__dfxtp_1
X_8102_ _7972_/B _8102_/B VGND VGND VPWR VPWR _8102_/X sky130_fd_sc_hd__and2b_1
X_6363_ _6363_/A _6363_/B VGND VGND VPWR VPWR _6414_/B sky130_fd_sc_hd__xnor2_1
X_9082_ _9224_/CLK _9082_/D VGND VGND VPWR VPWR _9082_/Q sky130_fd_sc_hd__dfxtp_1
X_5314_ _5314_/A VGND VGND VPWR VPWR _5315_/A sky130_fd_sc_hd__clkbuf_2
X_6294_ _6294_/A VGND VGND VPWR VPWR _6294_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8033_ _8033_/A _8033_/B VGND VGND VPWR VPWR _8116_/A sky130_fd_sc_hd__xor2_1
X_5245_ _5245_/A VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5176_ _5129_/X _5581_/A _5168_/X _5174_/Y _5175_/X VGND VGND VPWR VPWR _5176_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8935_ _8935_/A _8935_/B VGND VGND VPWR VPWR _8936_/B sky130_fd_sc_hd__and2_1
XFILLER_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8866_ _8866_/A _8866_/B VGND VGND VPWR VPWR _8868_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8797_ _8797_/A _8862_/A VGND VGND VPWR VPWR _8800_/A sky130_fd_sc_hd__xnor2_1
X_7817_ _7817_/A _7817_/B VGND VGND VPWR VPWR _7834_/A sky130_fd_sc_hd__or2_1
X_7748_ _7748_/A VGND VGND VPWR VPWR _8150_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_12_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7679_ _8867_/B VGND VGND VPWR VPWR _8816_/B sky130_fd_sc_hd__buf_2
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _9127_/Q _9119_/Q VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__and2_1
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6981_ _7078_/A _7078_/B VGND VGND VPWR VPWR _7106_/A sky130_fd_sc_hd__xnor2_1
X_8720_ _8720_/A _8720_/B VGND VGND VPWR VPWR _8887_/A sky130_fd_sc_hd__and2_2
X_5932_ _5929_/X _5930_/Y _5932_/B1 _5898_/X VGND VGND VPWR VPWR _5932_/X sky130_fd_sc_hd__a211o_1
XFILLER_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8651_ _8580_/Y _8579_/A _8578_/X VGND VGND VPWR VPWR _8772_/A sky130_fd_sc_hd__o21ai_1
X_5863_ _5863_/A _5863_/B _5863_/C VGND VGND VPWR VPWR _5898_/B sky130_fd_sc_hd__or3_1
X_7602_ _7602_/A _7849_/B VGND VGND VPWR VPWR _7606_/A sky130_fd_sc_hd__nand2_1
X_8582_ _8582_/A _8582_/B VGND VGND VPWR VPWR _9100_/D sky130_fd_sc_hd__xor2_1
X_4814_ _9124_/Q _9116_/Q VGND VGND VPWR VPWR _4815_/B sky130_fd_sc_hd__or2_1
X_5794_ _6885_/A VGND VGND VPWR VPWR _5908_/B sky130_fd_sc_hd__buf_2
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4745_ _4897_/A VGND VGND VPWR VPWR _5653_/B sky130_fd_sc_hd__buf_2
X_7533_ _7533_/A _7533_/B _7532_/Y VGND VGND VPWR VPWR _7535_/A sky130_fd_sc_hd__nor3b_1
X_7464_ _8093_/A _8268_/A VGND VGND VPWR VPWR _7470_/A sky130_fd_sc_hd__nand2_1
X_4676_ _4676_/A _4676_/B _4676_/C _4676_/D VGND VGND VPWR VPWR _4677_/C sky130_fd_sc_hd__or4_1
X_6415_ _8086_/A VGND VGND VPWR VPWR _8587_/A sky130_fd_sc_hd__clkbuf_2
X_9203_ _9219_/CLK _9203_/D VGND VGND VPWR VPWR _9203_/Q sky130_fd_sc_hd__dfxtp_2
X_7395_ _7394_/A _7394_/B _7393_/Y VGND VGND VPWR VPWR _7396_/B sky130_fd_sc_hd__o21ba_1
X_9134_ _9213_/CLK _9134_/D VGND VGND VPWR VPWR _9134_/Q sky130_fd_sc_hd__dfxtp_1
X_6346_ _6347_/B _6347_/C _6347_/A VGND VGND VPWR VPWR _6350_/A sky130_fd_sc_hd__a21o_1
X_9065_ _9065_/A _9065_/B VGND VGND VPWR VPWR _9161_/D sky130_fd_sc_hd__xor2_1
XFILLER_102_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8016_ _8016_/A _8016_/B VGND VGND VPWR VPWR _8018_/C sky130_fd_sc_hd__xnor2_1
X_6277_ _6927_/D VGND VGND VPWR VPWR _8243_/A sky130_fd_sc_hd__clkbuf_4
X_5228_ _5213_/X _5485_/A _5225_/X _5226_/Y _5227_/X VGND VGND VPWR VPWR _5228_/X
+ sky130_fd_sc_hd__a221o_1
X_5159_ _5138_/X _5430_/A _5153_/X _5157_/Y _5158_/X VGND VGND VPWR VPWR _5159_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8918_ _8918_/A _8963_/B VGND VGND VPWR VPWR _8920_/A sky130_fd_sc_hd__nor2_1
X_8849_ _8849_/A _8906_/A VGND VGND VPWR VPWR _8852_/A sky130_fd_sc_hd__xnor2_1
XFILLER_72_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6200_ _7610_/B VGND VGND VPWR VPWR _8156_/B sky130_fd_sc_hd__clkbuf_4
X_7180_ _7182_/A _7182_/B VGND VGND VPWR VPWR _7552_/A sky130_fd_sc_hd__xor2_2
X_6131_ _6131_/A VGND VGND VPWR VPWR _6132_/A sky130_fd_sc_hd__inv_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6702_/B VGND VGND VPWR VPWR _6925_/A sky130_fd_sc_hd__buf_2
XFILLER_58_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5013_ _5135_/A _5012_/Y _4926_/X VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__o21a_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6964_ _7923_/D VGND VGND VPWR VPWR _8175_/D sky130_fd_sc_hd__buf_2
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6895_ _7506_/A _7116_/D _7254_/D _5818_/X VGND VGND VPWR VPWR _6896_/B sky130_fd_sc_hd__a22oi_1
X_8703_ _8703_/A _8703_/B VGND VGND VPWR VPWR _8761_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5915_ _5915_/A _5915_/B _5915_/C VGND VGND VPWR VPWR _5918_/B sky130_fd_sc_hd__nand3_1
X_8634_ _8639_/A _8981_/B _8537_/A _8633_/X VGND VGND VPWR VPWR _8634_/Y sky130_fd_sc_hd__a31oi_1
X_5846_ _6660_/A _5922_/A VGND VGND VPWR VPWR _5847_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8565_ _8565_/A _8565_/B _8564_/Y VGND VGND VPWR VPWR _8567_/A sky130_fd_sc_hd__nor3b_1
X_5777_ _4587_/X _5776_/X _4870_/S VGND VGND VPWR VPWR _5777_/Y sky130_fd_sc_hd__o21ai_1
X_7516_ _7516_/A _7516_/B _7658_/A VGND VGND VPWR VPWR _7658_/B sky130_fd_sc_hd__nor3_2
X_8496_ _8496_/A _8496_/B VGND VGND VPWR VPWR _8498_/C sky130_fd_sc_hd__nor2_1
X_4728_ _9105_/Q VGND VGND VPWR VPWR _5736_/S sky130_fd_sc_hd__inv_2
X_7447_ _7447_/A _7447_/B _7447_/C VGND VGND VPWR VPWR _7447_/X sky130_fd_sc_hd__and3_1
X_4659_ _4659_/A VGND VGND VPWR VPWR _4660_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7378_ _7375_/X _7376_/Y _7377_/C _7377_/Y VGND VGND VPWR VPWR _7378_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_88_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9117_ _9218_/CLK hold18/X VGND VGND VPWR VPWR _9117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6329_ _6329_/A _6329_/B VGND VGND VPWR VPWR _6433_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9048_ _9022_/A _9022_/B _9040_/A _9047_/X VGND VGND VPWR VPWR _9049_/B sky130_fd_sc_hd__o31ai_2
XFILLER_57_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5700_ _5189_/X _4812_/X _5699_/X VGND VGND VPWR VPWR _9147_/D sky130_fd_sc_hd__o21ai_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6680_ _6680_/A _6680_/B _7327_/A _7042_/C VGND VGND VPWR VPWR _6805_/A sky130_fd_sc_hd__and4_1
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5631_ _5606_/X _5510_/X _5511_/X _5629_/X _5630_/X VGND VGND VPWR VPWR _9144_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8350_ _8521_/A _8351_/B _8348_/Y _8349_/X VGND VGND VPWR VPWR _8352_/A sky130_fd_sc_hd__o2bb2a_1
X_5562_ _5141_/A _5634_/A _5561_/X _5219_/A VGND VGND VPWR VPWR _5562_/X sky130_fd_sc_hd__a211o_1
X_8281_ _8498_/A _8846_/B VGND VGND VPWR VPWR _8282_/B sky130_fd_sc_hd__nand2_1
X_7301_ _7301_/A _7301_/B VGND VGND VPWR VPWR _7302_/B sky130_fd_sc_hd__and2_1
X_7232_ _7233_/A _7233_/B VGND VGND VPWR VPWR _7234_/A sky130_fd_sc_hd__or2_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5493_ _5165_/X _5206_/A _5491_/X _5492_/Y _5380_/X VGND VGND VPWR VPWR _5493_/X
+ sky130_fd_sc_hd__a221o_1
X_7163_ _7212_/B _7212_/C VGND VGND VPWR VPWR _7164_/B sky130_fd_sc_hd__nand2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6107_/X _6108_/X _6875_/A _8349_/A VGND VGND VPWR VPWR _6294_/A sky130_fd_sc_hd__o211a_2
X_7094_ _7094_/A _7094_/B VGND VGND VPWR VPWR _7097_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6045_ _6221_/A _6044_/C _6047_/B _6000_/A VGND VGND VPWR VPWR _6047_/D sky130_fd_sc_hd__o2bb2a_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7996_ _7997_/A _7997_/B VGND VGND VPWR VPWR _8081_/A sky130_fd_sc_hd__or2_1
XFILLER_81_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6947_ _6945_/C _6945_/Y _6943_/X _7059_/B VGND VGND VPWR VPWR _6948_/B sky130_fd_sc_hd__a211oi_1
XFILLER_22_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6878_ _6878_/A _6878_/B VGND VGND VPWR VPWR _6879_/C sky130_fd_sc_hd__and2_1
X_8617_ _8548_/A _8548_/B _8616_/X VGND VGND VPWR VPWR _8619_/B sky130_fd_sc_hd__a21oi_1
X_5829_ _6885_/A VGND VGND VPWR VPWR _6998_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8548_ _8548_/A _8548_/B VGND VGND VPWR VPWR _8551_/A sky130_fd_sc_hd__xnor2_1
X_8479_ _8480_/A _8480_/B VGND VGND VPWR VPWR _8479_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7850_ _7850_/A _7850_/B VGND VGND VPWR VPWR _7859_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6801_ _6801_/A _6801_/B VGND VGND VPWR VPWR _6802_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7781_ _7660_/A _7660_/B _7780_/X VGND VGND VPWR VPWR _7899_/B sky130_fd_sc_hd__a21o_1
X_4993_ _4994_/B _4993_/B VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__and2b_1
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6732_ _6853_/A _6732_/B VGND VGND VPWR VPWR _6734_/B sky130_fd_sc_hd__nor2_1
X_6663_ _6998_/A _6998_/B _6663_/C _7254_/D VGND VGND VPWR VPWR _6664_/B sky130_fd_sc_hd__and4_1
X_8402_ _8305_/B _8307_/Y _8399_/X _8494_/A VGND VGND VPWR VPWR _8494_/B sky130_fd_sc_hd__o211ai_4
X_5614_ _5424_/X _5136_/X _4558_/A VGND VGND VPWR VPWR _5614_/Y sky130_fd_sc_hd__a21oi_1
X_6594_ _6894_/A _7006_/B _6663_/C _7131_/C VGND VGND VPWR VPWR _6596_/A sky130_fd_sc_hd__and4_1
X_8333_ _8333_/A VGND VGND VPWR VPWR _8333_/Y sky130_fd_sc_hd__inv_2
X_5545_ _5245_/A _5170_/X _5543_/X _5544_/Y _5173_/X VGND VGND VPWR VPWR _5545_/X
+ sky130_fd_sc_hd__a221o_1
X_8264_ _8264_/A VGND VGND VPWR VPWR _8266_/B sky130_fd_sc_hd__inv_2
X_5476_ _5287_/A _5475_/X _5670_/S VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8195_ _8195_/A _8301_/B VGND VGND VPWR VPWR _8196_/B sky130_fd_sc_hd__xnor2_1
X_7215_ _7215_/A VGND VGND VPWR VPWR _7215_/Y sky130_fd_sc_hd__inv_2
X_7146_ _7146_/A _7730_/B VGND VGND VPWR VPWR _7150_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _7077_/A _7077_/B _7079_/B VGND VGND VPWR VPWR _7088_/A sky130_fd_sc_hd__or3_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6028_ _6022_/A _7348_/A _7347_/A _5985_/A VGND VGND VPWR VPWR _6029_/B sky130_fd_sc_hd__a22oi_1
XFILLER_27_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7979_ _7976_/Y _8064_/A _7978_/X _7860_/B VGND VGND VPWR VPWR _7981_/A sky130_fd_sc_hd__a211o_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5330_ _5206_/A _5329_/X _5354_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
X_5261_ _5160_/X _5507_/A _4599_/A VGND VGND VPWR VPWR _5261_/Y sky130_fd_sc_hd__a21oi_1
X_7000_ _6530_/B _7116_/D _7988_/B _6886_/A VGND VGND VPWR VPWR _7000_/Y sky130_fd_sc_hd__a22oi_1
X_5192_ _9087_/Q VGND VGND VPWR VPWR _5205_/A sky130_fd_sc_hd__buf_2
X_8951_ _8951_/A _8951_/B VGND VGND VPWR VPWR _8952_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7902_ _7902_/A _7902_/B VGND VGND VPWR VPWR _7903_/C sky130_fd_sc_hd__xnor2_1
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8882_ _8775_/B _8880_/Y _8881_/X VGND VGND VPWR VPWR _8884_/B sky130_fd_sc_hd__a21o_1
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7833_ _7834_/A _7834_/B VGND VGND VPWR VPWR _7837_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7764_ _7764_/A _7764_/B VGND VGND VPWR VPWR _7772_/B sky130_fd_sc_hd__and2_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6715_ _6814_/A _6814_/B _6814_/C VGND VGND VPWR VPWR _6715_/X sky130_fd_sc_hd__or3_1
X_4976_ _4932_/X _4933_/Y _5305_/S VGND VGND VPWR VPWR _4976_/X sky130_fd_sc_hd__a21o_1
X_7695_ _7696_/C _7571_/A _7693_/Y _7694_/X VGND VGND VPWR VPWR _7697_/A sky130_fd_sc_hd__o2bb2a_1
X_6646_ _6646_/A _6646_/B VGND VGND VPWR VPWR _6655_/C sky130_fd_sc_hd__xor2_2
X_6577_ _6502_/B _6504_/B _6502_/A VGND VGND VPWR VPWR _6578_/B sky130_fd_sc_hd__o21ba_1
X_8316_ _8181_/B _8316_/B VGND VGND VPWR VPWR _8316_/X sky130_fd_sc_hd__and2b_1
X_5528_ _5402_/A _5527_/X _5575_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8247_ _8607_/D VGND VGND VPWR VPWR _8664_/C sky130_fd_sc_hd__clkbuf_2
X_5459_ _5433_/X _5365_/X _5366_/X _5457_/X _5458_/X VGND VGND VPWR VPWR _9137_/D
+ sky130_fd_sc_hd__o221a_2
X_8178_ _8415_/A _8597_/B VGND VGND VPWR VPWR _8179_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7129_ _7129_/A _7129_/B VGND VGND VPWR VPWR _7133_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4830_ _4939_/A _4957_/A VGND VGND VPWR VPWR _4830_/X sky130_fd_sc_hd__or2b_4
X_4761_ _4837_/A _4762_/A VGND VGND VPWR VPWR _4929_/A sky130_fd_sc_hd__and2_1
XFILLER_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7480_ _7847_/D VGND VGND VPWR VPWR _8290_/A sky130_fd_sc_hd__clkbuf_4
X_6500_ _7293_/B _6500_/B _6759_/C _6927_/D VGND VGND VPWR VPWR _6502_/A sky130_fd_sc_hd__and4_1
X_4692_ _4828_/A VGND VGND VPWR VPWR _4842_/A sky130_fd_sc_hd__clkbuf_2
X_6431_ _6488_/A _6431_/B VGND VGND VPWR VPWR _6432_/B sky130_fd_sc_hd__xnor2_1
X_9150_ _9199_/CLK _9150_/D VGND VGND VPWR VPWR _9150_/Q sky130_fd_sc_hd__dfxtp_1
X_6362_ _6362_/A _6362_/B VGND VGND VPWR VPWR _6363_/B sky130_fd_sc_hd__nor2_1
X_8101_ _8100_/A _8100_/B _8100_/C VGND VGND VPWR VPWR _8203_/A sky130_fd_sc_hd__a21o_2
X_5313_ _5313_/A VGND VGND VPWR VPWR _5314_/A sky130_fd_sc_hd__clkbuf_2
X_9081_ _9214_/CLK _9081_/D VGND VGND VPWR VPWR _9081_/Q sky130_fd_sc_hd__dfxtp_1
X_6293_ _6293_/A _6378_/B VGND VGND VPWR VPWR _6380_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8032_ _8032_/A _8867_/B VGND VGND VPWR VPWR _8033_/B sky130_fd_sc_hd__nand2_1
X_5244_ _5244_/A VGND VGND VPWR VPWR _5245_/A sky130_fd_sc_hd__clkbuf_2
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5175_ _5175_/A VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8934_ _8935_/A _8935_/B VGND VGND VPWR VPWR _8936_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8865_ _8865_/A _8865_/B _8865_/C VGND VGND VPWR VPWR _8866_/B sky130_fd_sc_hd__and3_1
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7816_ _7816_/A _7816_/B VGND VGND VPWR VPWR _7817_/B sky130_fd_sc_hd__and2_1
X_8796_ _8734_/A _8736_/B _8734_/B VGND VGND VPWR VPWR _8862_/A sky130_fd_sc_hd__o21ba_1
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7747_ _8137_/A VGND VGND VPWR VPWR _7747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4959_ _5382_/A _4956_/X _4957_/Y _4958_/X VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__o22a_1
X_7678_ _7796_/B _7678_/B VGND VGND VPWR VPWR _9091_/D sky130_fd_sc_hd__nor2_1
X_6629_ _7962_/B VGND VGND VPWR VPWR _8519_/A sky130_fd_sc_hd__buf_4
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6980_ _7077_/A _6980_/B VGND VGND VPWR VPWR _7078_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5931_ _5931_/A1 _5898_/X _5929_/X _5930_/Y VGND VGND VPWR VPWR _6000_/A sky130_fd_sc_hd__o211ai_4
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8650_ _8429_/B _8510_/Y _8582_/A _8427_/B _8512_/A VGND VGND VPWR VPWR _8652_/B
+ sky130_fd_sc_hd__a2111o_1
X_5862_ _5863_/B _5863_/C _5863_/A VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__o21a_1
X_7601_ _7601_/A _7601_/B VGND VGND VPWR VPWR _7616_/B sky130_fd_sc_hd__nand2_1
X_8581_ _8512_/A _8512_/B _8580_/Y VGND VGND VPWR VPWR _8582_/B sky130_fd_sc_hd__o21ba_1
X_4813_ _9124_/Q _9116_/Q VGND VGND VPWR VPWR _4901_/A sky130_fd_sc_hd__nand2_1
X_5793_ _9197_/Q VGND VGND VPWR VPWR _6885_/A sky130_fd_sc_hd__clkbuf_2
X_4744_ _5510_/A _4966_/B _4743_/X VGND VGND VPWR VPWR _4744_/Y sky130_fd_sc_hd__o21ai_1
X_7532_ _7298_/A _7298_/B _7302_/B VGND VGND VPWR VPWR _7532_/Y sky130_fd_sc_hd__a21oi_1
X_7463_ _8050_/A VGND VGND VPWR VPWR _8268_/A sky130_fd_sc_hd__buf_2
X_4675_ _5364_/A _5460_/A _5271_/A _4675_/D VGND VGND VPWR VPWR _4676_/D sky130_fd_sc_hd__or4_1
X_9202_ _9216_/CLK _9202_/D VGND VGND VPWR VPWR _9202_/Q sky130_fd_sc_hd__dfxtp_2
X_6414_ _6365_/B _6414_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2b_1
X_7394_ _7394_/A _7394_/B _7393_/Y VGND VGND VPWR VPWR _7396_/A sky130_fd_sc_hd__nor3b_1
X_9133_ _9213_/CLK _9133_/D VGND VGND VPWR VPWR _9133_/Q sky130_fd_sc_hd__dfxtp_1
X_6345_ _6345_/A _6387_/B VGND VGND VPWR VPWR _6347_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6276_ _7042_/D VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_9064_ _9064_/A _9064_/B VGND VGND VPWR VPWR _9068_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8015_ _8122_/A _8015_/B VGND VGND VPWR VPWR _8016_/B sky130_fd_sc_hd__xnor2_1
X_5227_ _5227_/A VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5158_ _5158_/A VGND VGND VPWR VPWR _5158_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5089_ _5187_/A _4932_/X _5067_/X _9109_/Q VGND VGND VPWR VPWR _5089_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8917_ _8914_/Y _8917_/B VGND VGND VPWR VPWR _8963_/B sky130_fd_sc_hd__and2b_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8848_ _8793_/A _8795_/B _8793_/B VGND VGND VPWR VPWR _8906_/A sky130_fd_sc_hd__o21ba_1
XFILLER_72_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8779_ _8780_/A _8780_/B _8887_/A VGND VGND VPWR VPWR _8781_/A sky130_fd_sc_hd__a21oi_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6130_ _6125_/A _6126_/X _6125_/B VGND VGND VPWR VPWR _6218_/B sky130_fd_sc_hd__a21o_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6702_/A VGND VGND VPWR VPWR _6572_/B sky130_fd_sc_hd__clkbuf_2
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5003_/X _4929_/B _5011_/Y VGND VGND VPWR VPWR _5012_/Y sky130_fd_sc_hd__a21oi_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6963_ _7419_/D VGND VGND VPWR VPWR _7923_/D sky130_fd_sc_hd__clkbuf_2
X_6894_ _6894_/A _7119_/B _7347_/B _7348_/B VGND VGND VPWR VPWR _6896_/A sky130_fd_sc_hd__and4_1
XFILLER_81_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8702_ _8703_/A _8703_/B VGND VGND VPWR VPWR _8704_/A sky130_fd_sc_hd__and2_1
X_5914_ _5915_/A _5915_/B _5915_/C VGND VGND VPWR VPWR _5918_/A sky130_fd_sc_hd__a21o_1
X_8633_ _8535_/B _8633_/B VGND VGND VPWR VPWR _8633_/X sky130_fd_sc_hd__and2b_1
XFILLER_22_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5845_ _9198_/Q VGND VGND VPWR VPWR _6660_/A sky130_fd_sc_hd__buf_2
XFILLER_61_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8564_ _8568_/A _8981_/B _8460_/A _8563_/X VGND VGND VPWR VPWR _8564_/Y sky130_fd_sc_hd__a31oi_1
X_5776_ _5314_/A _4573_/A _4580_/X _5244_/A _4566_/X VGND VGND VPWR VPWR _5776_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7515_ _7514_/A _7514_/B _7514_/C VGND VGND VPWR VPWR _7658_/A sky130_fd_sc_hd__o21a_1
X_8495_ _8494_/A _8494_/B _8494_/C VGND VGND VPWR VPWR _8496_/B sky130_fd_sc_hd__a21oi_2
X_4727_ _4720_/X _4725_/Y _4726_/X _4966_/B VGND VGND VPWR VPWR _4727_/X sky130_fd_sc_hd__o2bb2a_1
X_7446_ _7446_/A _7446_/B VGND VGND VPWR VPWR _7447_/C sky130_fd_sc_hd__nand2_1
X_4658_ _4658_/A VGND VGND VPWR VPWR _4659_/A sky130_fd_sc_hd__clkbuf_2
X_9116_ _9116_/CLK hold4/X VGND VGND VPWR VPWR _9116_/Q sky130_fd_sc_hd__dfxtp_2
X_7377_ _7377_/A _7377_/B _7377_/C VGND VGND VPWR VPWR _7377_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4589_ _9097_/Q VGND VGND VPWR VPWR _4839_/A sky130_fd_sc_hd__clkbuf_2
X_6328_ _6328_/A _6328_/B VGND VGND VPWR VPWR _6433_/A sky130_fd_sc_hd__xnor2_4
XFILLER_103_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9047_ _9038_/Y _9037_/A _9036_/X VGND VGND VPWR VPWR _9047_/X sky130_fd_sc_hd__o21a_1
X_6259_ _6259_/A _6259_/B VGND VGND VPWR VPWR _6351_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5630_ _5630_/A _5653_/B VGND VGND VPWR VPWR _5630_/X sky130_fd_sc_hd__or2_1
X_5561_ _4570_/A _5607_/A _5559_/Y _5560_/X _5007_/A VGND VGND VPWR VPWR _5561_/X
+ sky130_fd_sc_hd__o221a_1
X_8280_ _8597_/B VGND VGND VPWR VPWR _8846_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5492_ _5247_/X _5656_/A _5378_/X VGND VGND VPWR VPWR _5492_/Y sky130_fd_sc_hd__a21oi_1
X_7300_ _7301_/A _7301_/B VGND VGND VPWR VPWR _7302_/A sky130_fd_sc_hd__nor2_1
X_7231_ _7231_/A _7342_/C VGND VGND VPWR VPWR _7233_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7162_ _7161_/A _7161_/B _7161_/C VGND VGND VPWR VPWR _7212_/C sky130_fd_sc_hd__a21o_2
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6113_ _8154_/A VGND VGND VPWR VPWR _8349_/A sky130_fd_sc_hd__buf_4
XFILLER_86_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7187_/B _7093_/B _7694_/C _7694_/D VGND VGND VPWR VPWR _7094_/B sky130_fd_sc_hd__and4_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6044_ _6000_/A _6047_/B _6044_/C _6221_/A VGND VGND VPWR VPWR _6131_/A sky130_fd_sc_hd__and4bb_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7995_ _7995_/A _8083_/A VGND VGND VPWR VPWR _7997_/B sky130_fd_sc_hd__xor2_1
XFILLER_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6946_ _6943_/X _7059_/B _6945_/C _6945_/Y VGND VGND VPWR VPWR _6948_/A sky130_fd_sc_hd__o211a_1
XFILLER_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6877_ _6877_/A _6877_/B VGND VGND VPWR VPWR _6878_/B sky130_fd_sc_hd__or2_1
X_8616_ _8547_/A _8616_/B VGND VGND VPWR VPWR _8616_/X sky130_fd_sc_hd__and2b_1
X_5828_ _6974_/B VGND VGND VPWR VPWR _7293_/B sky130_fd_sc_hd__clkbuf_2
X_8547_ _8547_/A _8616_/B VGND VGND VPWR VPWR _8548_/B sky130_fd_sc_hd__xnor2_1
X_5759_ _5534_/X _5606_/X _5758_/X _4999_/X VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__o31a_1
X_8478_ _8478_/A _8478_/B VGND VGND VPWR VPWR _8480_/B sky130_fd_sc_hd__nand2_1
X_7429_ _7429_/A _7429_/B VGND VGND VPWR VPWR _7445_/A sky130_fd_sc_hd__or2_1
XFILLER_103_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6800_ _5985_/D _7327_/B _7330_/A _6172_/A VGND VGND VPWR VPWR _6801_/B sky130_fd_sc_hd__a22oi_1
X_7780_ _7659_/B _7780_/B VGND VGND VPWR VPWR _7780_/X sky130_fd_sc_hd__and2b_1
X_4992_ _4992_/A _5033_/A VGND VGND VPWR VPWR _4993_/B sky130_fd_sc_hd__or2_1
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6731_ _6730_/B _6730_/C _6730_/A VGND VGND VPWR VPWR _6732_/B sky130_fd_sc_hd__a21oi_1
X_6662_ _6530_/B _7129_/B _7254_/D _6886_/A VGND VGND VPWR VPWR _6664_/A sky130_fd_sc_hd__a22oi_2
XFILLER_31_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8401_ _8399_/X _8494_/A _8305_/B _8307_/Y VGND VGND VPWR VPWR _8403_/B sky130_fd_sc_hd__a211o_1
X_5613_ _5393_/A _5258_/X _5611_/X _5612_/Y _5410_/X VGND VGND VPWR VPWR _5613_/X
+ sky130_fd_sc_hd__a221o_1
X_6593_ _6593_/A _6886_/B VGND VGND VPWR VPWR _6597_/A sky130_fd_sc_hd__nand2_1
X_8332_ _8510_/A _8332_/B VGND VGND VPWR VPWR _8335_/A sky130_fd_sc_hd__and2b_1
X_5544_ _5394_/X _5132_/X _5414_/X VGND VGND VPWR VPWR _5544_/Y sky130_fd_sc_hd__a21oi_1
X_8263_ _8365_/A _8263_/B VGND VGND VPWR VPWR _8264_/A sky130_fd_sc_hd__nand2_1
X_5475_ _5245_/A _5474_/Y _5572_/S VGND VGND VPWR VPWR _5475_/X sky130_fd_sc_hd__mux2_1
X_8194_ _8194_/A _8299_/B VGND VGND VPWR VPWR _8301_/B sky130_fd_sc_hd__nor2_1
X_7214_ _7212_/C _7212_/Y _7210_/X _7211_/Y VGND VGND VPWR VPWR _7394_/A sky130_fd_sc_hd__a211oi_4
X_7145_ _7145_/A _7025_/B VGND VGND VPWR VPWR _7161_/B sky130_fd_sc_hd__or2b_1
XFILLER_59_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _7076_/A _7076_/B VGND VGND VPWR VPWR _7104_/B sky130_fd_sc_hd__or2_1
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6027_ _9200_/Q VGND VGND VPWR VPWR _7347_/A sky130_fd_sc_hd__clkbuf_2
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7978_ _7857_/B _7978_/B VGND VGND VPWR VPWR _7978_/X sky130_fd_sc_hd__and2b_1
X_6929_ _6929_/A _6929_/B VGND VGND VPWR VPWR _6930_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5260_ _9077_/Q VGND VGND VPWR VPWR _5507_/A sky130_fd_sc_hd__clkbuf_4
X_5191_ _4737_/X _5122_/X _5186_/X _5190_/Y _4739_/A VGND VGND VPWR VPWR _5191_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_95_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8950_ _8951_/A _8951_/B VGND VGND VPWR VPWR _8952_/A sky130_fd_sc_hd__or2_1
XFILLER_56_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7901_ _7901_/A _8013_/A VGND VGND VPWR VPWR _7902_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8881_ _8769_/A _8826_/A _8825_/Y VGND VGND VPWR VPWR _8881_/X sky130_fd_sc_hd__o21a_1
X_7832_ _7832_/A _7832_/B VGND VGND VPWR VPWR _7834_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7763_ _7763_/A _7845_/A VGND VGND VPWR VPWR _7865_/A sky130_fd_sc_hd__xnor2_4
X_4975_ _5739_/S VGND VGND VPWR VPWR _5305_/S sky130_fd_sc_hd__buf_2
X_6714_ _6814_/B _6814_/C _6814_/A VGND VGND VPWR VPWR _6714_/Y sky130_fd_sc_hd__o21ai_2
X_7694_ _7694_/A _7694_/B _7694_/C _7694_/D VGND VGND VPWR VPWR _7694_/X sky130_fd_sc_hd__and4_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6645_ _6656_/A _6656_/B VGND VGND VPWR VPWR _6646_/B sky130_fd_sc_hd__xnor2_2
X_6576_ _6576_/A _6576_/B VGND VGND VPWR VPWR _6693_/B sky130_fd_sc_hd__xnor2_2
X_8315_ _8171_/X _8210_/B _8312_/Y _8313_/X VGND VGND VPWR VPWR _8421_/A sky130_fd_sc_hd__a211oi_2
X_5527_ _5364_/A _5526_/X _5527_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
X_8246_ _8154_/X _8522_/A _8245_/Y VGND VGND VPWR VPWR _8249_/A sky130_fd_sc_hd__a21oi_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5458_ _9075_/Q _5482_/B VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__or2_1
X_8177_ _8177_/A VGND VGND VPWR VPWR _8415_/A sky130_fd_sc_hd__clkbuf_2
X_5389_ _5389_/A VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__clkbuf_2
X_7128_ _7021_/A _7020_/A _7020_/B VGND VGND VPWR VPWR _7219_/A sky130_fd_sc_hd__o21ba_1
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7059_ _7059_/A _7059_/B VGND VGND VPWR VPWR _7060_/B sky130_fd_sc_hd__nor2_2
XFILLER_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4760_ _4852_/A _4866_/A VGND VGND VPWR VPWR _4760_/X sky130_fd_sc_hd__or2_2
X_4691_ _4691_/A _4691_/B VGND VGND VPWR VPWR _4828_/A sky130_fd_sc_hd__nand2_1
X_6430_ _6430_/A _6430_/B VGND VGND VPWR VPWR _6431_/B sky130_fd_sc_hd__xnor2_2
X_6361_ _7081_/A _6361_/B _6361_/C _6361_/D VGND VGND VPWR VPWR _6362_/B sky130_fd_sc_hd__and4_1
X_8100_ _8100_/A _8100_/B _8100_/C VGND VGND VPWR VPWR _8100_/Y sky130_fd_sc_hd__nand3_2
X_5312_ _5287_/X _5202_/X _5204_/X _5310_/X _5311_/X VGND VGND VPWR VPWR _9132_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9080_ _9214_/CLK _9080_/D VGND VGND VPWR VPWR _9080_/Q sky130_fd_sc_hd__dfxtp_1
X_6292_ _6292_/A _6292_/B _6378_/A VGND VGND VPWR VPWR _6378_/B sky130_fd_sc_hd__nand3_1
X_8031_ _8031_/A _8031_/B VGND VGND VPWR VPWR _8033_/A sky130_fd_sc_hd__nor2_1
X_5243_ _5200_/X _5202_/X _5204_/X _5241_/X _5242_/X VGND VGND VPWR VPWR _9130_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_102_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5174_ _5170_/X _5485_/A _5173_/X VGND VGND VPWR VPWR _5174_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8933_ _8989_/A _8933_/B VGND VGND VPWR VPWR _8935_/B sky130_fd_sc_hd__and2_1
X_8864_ _8865_/A _8865_/B _8865_/C VGND VGND VPWR VPWR _8866_/A sky130_fd_sc_hd__a21oi_1
XFILLER_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7815_ _7816_/A _7816_/B VGND VGND VPWR VPWR _7817_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8795_ _8795_/A _8795_/B VGND VGND VPWR VPWR _8797_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7746_ _7746_/A _7746_/B VGND VGND VPWR VPWR _7779_/A sky130_fd_sc_hd__nor2_2
X_4958_ _4957_/A _4957_/B _5732_/S VGND VGND VPWR VPWR _4958_/X sky130_fd_sc_hd__a21o_1
X_7677_ _7677_/A _7677_/B _7677_/C VGND VGND VPWR VPWR _7678_/B sky130_fd_sc_hd__and3_1
X_4889_ _4889_/A VGND VGND VPWR VPWR _4889_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6628_ _8542_/A VGND VGND VPWR VPWR _8780_/A sky130_fd_sc_hd__buf_4
X_6559_ _6478_/B _6480_/X _6558_/X VGND VGND VPWR VPWR _6649_/A sky130_fd_sc_hd__a21oi_2
XFILLER_105_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8229_ _8229_/A _8229_/B _8229_/C VGND VGND VPWR VPWR _8333_/A sky130_fd_sc_hd__and3_1
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5930_ _5930_/A _5930_/B _5930_/C VGND VGND VPWR VPWR _5930_/Y sky130_fd_sc_hd__nand3_2
X_7600_ _7600_/A _7493_/B VGND VGND VPWR VPWR _7616_/A sky130_fd_sc_hd__or2b_1
XFILLER_61_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5861_ _5861_/A _5861_/B VGND VGND VPWR VPWR _5863_/A sky130_fd_sc_hd__xor2_2
X_8580_ _8580_/A _8580_/B VGND VGND VPWR VPWR _8580_/Y sky130_fd_sc_hd__nor2_1
X_5792_ _6151_/A VGND VGND VPWR VPWR _5945_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4812_ _5785_/S VGND VGND VPWR VPWR _4812_/X sky130_fd_sc_hd__buf_2
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4743_ _4687_/X _4693_/Y _4741_/Y _4896_/A VGND VGND VPWR VPWR _4743_/X sky130_fd_sc_hd__a211o_1
X_7531_ _7531_/A _7804_/B VGND VGND VPWR VPWR _7536_/A sky130_fd_sc_hd__nand2_1
X_7462_ _7462_/A VGND VGND VPWR VPWR _8093_/A sky130_fd_sc_hd__clkbuf_2
X_9201_ _9208_/CLK _9201_/D VGND VGND VPWR VPWR _9201_/Q sky130_fd_sc_hd__dfxtp_4
X_6413_ _6483_/B VGND VGND VPWR VPWR _6413_/Y sky130_fd_sc_hd__inv_2
X_4674_ _5244_/A _5200_/A _4874_/S _5385_/A VGND VGND VPWR VPWR _4675_/D sky130_fd_sc_hd__or4_1
X_7393_ _7389_/A _8850_/B _7195_/A _7392_/X VGND VGND VPWR VPWR _7393_/Y sky130_fd_sc_hd__a31oi_1
X_9132_ _9214_/CLK _9132_/D VGND VGND VPWR VPWR _9132_/Q sky130_fd_sc_hd__dfxtp_1
X_6344_ _6344_/A _6411_/A VGND VGND VPWR VPWR _6387_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9063_ _5945_/A _7531_/A _7389_/A _7645_/A VGND VGND VPWR VPWR _9064_/B sky130_fd_sc_hd__a22oi_2
X_6275_ _6567_/B _6858_/A _7852_/A _7610_/B VGND VGND VPWR VPWR _6279_/A sky130_fd_sc_hd__and4_1
X_8014_ _7902_/A _7902_/B _8013_/X VGND VGND VPWR VPWR _8015_/B sky130_fd_sc_hd__a21bo_1
X_5226_ _4717_/S _5532_/A _4605_/A VGND VGND VPWR VPWR _5226_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5157_ _5154_/X _5316_/A _5156_/X VGND VGND VPWR VPWR _5157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5088_ _4932_/X _4998_/A _5041_/A _5695_/S VGND VGND VPWR VPWR _5088_/Y sky130_fd_sc_hd__a211oi_1
X_8916_ _8916_/A _8963_/A VGND VGND VPWR VPWR _8917_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8847_ _8847_/A _8847_/B VGND VGND VPWR VPWR _8849_/A sky130_fd_sc_hd__xnor2_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8778_ _8778_/A _8814_/A _8778_/C VGND VGND VPWR VPWR _8809_/A sky130_fd_sc_hd__or3_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7729_ _7729_/A _7729_/B VGND VGND VPWR VPWR _7731_/A sky130_fd_sc_hd__nor2_1
XANTENNA_60 _9130_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6223_/A _6223_/B _7037_/A _7148_/A VGND VGND VPWR VPWR _6068_/B sky130_fd_sc_hd__nand4_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5011_ _4947_/Y _5010_/X _5058_/A VGND VGND VPWR VPWR _5011_/Y sky130_fd_sc_hd__a21oi_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6962_ _9212_/Q VGND VGND VPWR VPWR _7419_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6893_ _7118_/A _7360_/A VGND VGND VPWR VPWR _6897_/A sky130_fd_sc_hd__nand2_1
X_8701_ _8701_/A _8701_/B VGND VGND VPWR VPWR _8703_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5913_ _5913_/A _5913_/B VGND VGND VPWR VPWR _5915_/C sky130_fd_sc_hd__xnor2_1
X_8632_ _8632_/A _8705_/A VGND VGND VPWR VPWR _8656_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5844_ _5844_/A _5844_/B VGND VGND VPWR VPWR _5847_/A sky130_fd_sc_hd__nor2_1
X_8563_ _8458_/B _8563_/B VGND VGND VPWR VPWR _8563_/X sky130_fd_sc_hd__and2b_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7514_ _7514_/A _7514_/B _7514_/C VGND VGND VPWR VPWR _7516_/B sky130_fd_sc_hd__nor3_1
X_5775_ _4889_/X _5774_/X _5628_/A VGND VGND VPWR VPWR _5775_/X sky130_fd_sc_hd__o21a_1
X_8494_ _8494_/A _8494_/B _8494_/C VGND VGND VPWR VPWR _8496_/A sky130_fd_sc_hd__and3_1
X_4726_ _5691_/S VGND VGND VPWR VPWR _4726_/X sky130_fd_sc_hd__clkbuf_2
X_7445_ _7445_/A _7445_/B VGND VGND VPWR VPWR _7446_/B sky130_fd_sc_hd__or2_1
X_4657_ _4780_/A _4776_/A VGND VGND VPWR VPWR _4658_/A sky130_fd_sc_hd__or2_1
X_7376_ _7518_/B _7518_/C _7518_/A VGND VGND VPWR VPWR _7376_/Y sky130_fd_sc_hd__a21oi_1
X_9115_ _9210_/CLK hold12/X VGND VGND VPWR VPWR _9115_/Q sky130_fd_sc_hd__dfxtp_4
X_6327_ _6327_/A _6327_/B VGND VGND VPWR VPWR _6328_/B sky130_fd_sc_hd__nor2_2
X_4588_ _4573_/X _4580_/X _4587_/X VGND VGND VPWR VPWR _4588_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9046_ _9046_/A _9046_/B VGND VGND VPWR VPWR _9049_/A sky130_fd_sc_hd__xnor2_2
X_6258_ _6258_/A _6258_/B VGND VGND VPWR VPWR _6259_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6189_ _7152_/C VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5209_ _9083_/Q VGND VGND VPWR VPWR _5210_/A sky130_fd_sc_hd__buf_2
XFILLER_84_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5560_ _4849_/A _5184_/A _5146_/A _5179_/A _4783_/X VGND VGND VPWR VPWR _5560_/X
+ sky130_fd_sc_hd__a221o_1
X_5491_ _5160_/X _5208_/A _5489_/X _5490_/Y _5410_/X VGND VGND VPWR VPWR _5491_/X
+ sky130_fd_sc_hd__a221o_1
X_7230_ _7230_/A _7230_/B VGND VGND VPWR VPWR _7342_/C sky130_fd_sc_hd__nor2_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7161_ _7161_/A _7161_/B _7161_/C VGND VGND VPWR VPWR _7212_/B sky130_fd_sc_hd__nand3_4
X_6112_ _6361_/C VGND VGND VPWR VPWR _8154_/A sky130_fd_sc_hd__clkbuf_2
X_7092_ _9212_/Q VGND VGND VPWR VPWR _7694_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _5997_/B _5999_/A _6040_/Y _6041_/X VGND VGND VPWR VPWR _6221_/A sky130_fd_sc_hd__a211o_2
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7994_ _7994_/A _8100_/A VGND VGND VPWR VPWR _8083_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6945_ _6945_/A _6945_/B _6945_/C VGND VGND VPWR VPWR _6945_/Y sky130_fd_sc_hd__nand3_1
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6876_ _6877_/A _6877_/B VGND VGND VPWR VPWR _6878_/A sky130_fd_sc_hd__nand2_1
X_8615_ _8672_/B _8615_/B VGND VGND VPWR VPWR _8619_/A sky130_fd_sc_hd__nand2_1
X_5827_ _5834_/A _5834_/B VGND VGND VPWR VPWR _5863_/B sky130_fd_sc_hd__and2_1
X_8546_ _8546_/A _8614_/B VGND VGND VPWR VPWR _8616_/B sky130_fd_sc_hd__nor2_1
X_5758_ _5433_/X _5509_/A _5757_/X _5712_/S VGND VGND VPWR VPWR _5758_/X sky130_fd_sc_hd__o31a_1
X_8477_ _8477_/A _8477_/B VGND VGND VPWR VPWR _8478_/B sky130_fd_sc_hd__or2_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4709_ _4698_/X _4708_/X _5727_/S VGND VGND VPWR VPWR _4709_/X sky130_fd_sc_hd__mux2_1
X_7428_ _7428_/A _7428_/B VGND VGND VPWR VPWR _7429_/B sky130_fd_sc_hd__and2_1
X_5689_ _5156_/A _5227_/A _5687_/X _5688_/Y VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7359_ _7359_/A _9184_/Q _7503_/C VGND VGND VPWR VPWR _7482_/A sky130_fd_sc_hd__and3_1
XFILLER_103_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9029_ _9029_/A _9029_/B _9029_/C VGND VGND VPWR VPWR _9031_/A sky130_fd_sc_hd__and3_1
XFILLER_1_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ _4991_/A _4991_/B VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__nor2_1
X_6730_ _6730_/A _6730_/B _6730_/C VGND VGND VPWR VPWR _6853_/A sky130_fd_sc_hd__and3_1
X_6661_ _9178_/Q VGND VGND VPWR VPWR _7254_/D sky130_fd_sc_hd__buf_2
XFILLER_31_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8400_ _8255_/B _8398_/X _8396_/Y _8397_/X VGND VGND VPWR VPWR _8494_/A sky130_fd_sc_hd__o211ai_4
X_6592_ _6592_/A _6592_/B VGND VGND VPWR VPWR _6659_/A sky130_fd_sc_hd__xnor2_1
X_5612_ _5138_/X _5420_/X _5158_/X VGND VGND VPWR VPWR _5612_/Y sky130_fd_sc_hd__a21oi_1
X_8331_ _8331_/A _8331_/B _8329_/Y VGND VGND VPWR VPWR _8332_/B sky130_fd_sc_hd__or3b_1
X_5543_ _5165_/X _5116_/A _5541_/X _5542_/Y _5380_/X VGND VGND VPWR VPWR _5543_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8262_ _7747_/X _8978_/B _8257_/C _8257_/B VGND VGND VPWR VPWR _8263_/B sky130_fd_sc_hd__a31o_1
X_5474_ _5394_/X _4966_/A _5473_/X VGND VGND VPWR VPWR _5474_/Y sky130_fd_sc_hd__o21ai_1
X_8193_ _8268_/A _8467_/A _8193_/C VGND VGND VPWR VPWR _8299_/B sky130_fd_sc_hd__and3_1
X_7213_ _7210_/X _7211_/Y _7212_/C _7212_/Y VGND VGND VPWR VPWR _7213_/X sky130_fd_sc_hd__o211a_1
X_7144_ _7047_/A _7047_/B _7143_/X VGND VGND VPWR VPWR _7164_/A sky130_fd_sc_hd__a21oi_2
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7075_/A _7174_/B _7075_/C VGND VGND VPWR VPWR _7172_/B sky130_fd_sc_hd__or3_1
XFILLER_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6026_ _9199_/Q VGND VGND VPWR VPWR _7348_/A sky130_fd_sc_hd__buf_2
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7977_ _7976_/A _7976_/B _7976_/C VGND VGND VPWR VPWR _8064_/A sky130_fd_sc_hd__a21o_2
XFILLER_54_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6928_ _7583_/B _6361_/C _7610_/B _6679_/A VGND VGND VPWR VPWR _6929_/B sky130_fd_sc_hd__a22oi_1
XFILLER_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6859_ _6859_/A _6859_/B _7822_/C _7822_/D VGND VGND VPWR VPWR _6861_/A sky130_fd_sc_hd__and4_1
XFILLER_80_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8529_ _8532_/D VGND VGND VPWR VPWR _8529_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5190_ _5187_/X _5189_/X _4737_/A VGND VGND VPWR VPWR _5190_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7900_ _7783_/A _7783_/B _7899_/X VGND VGND VPWR VPWR _8013_/A sky130_fd_sc_hd__a21oi_1
X_8880_ _8880_/A _8880_/B VGND VGND VPWR VPWR _8880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7831_ _7830_/A _7830_/B _7829_/X VGND VGND VPWR VPWR _7832_/B sky130_fd_sc_hd__o21bai_1
X_7762_ _7762_/A _7861_/A VGND VGND VPWR VPWR _7845_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4974_ _5236_/S _4969_/X _4972_/Y _4973_/X VGND VGND VPWR VPWR _4974_/X sky130_fd_sc_hd__a31o_1
X_7693_ _7696_/D VGND VGND VPWR VPWR _7693_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6713_ _6817_/A _6817_/B VGND VGND VPWR VPWR _6814_/A sky130_fd_sc_hd__xnor2_2
X_6644_ _6553_/A _6642_/X _6643_/Y VGND VGND VPWR VPWR _6656_/B sky130_fd_sc_hd__a21bo_1
X_6575_ _7419_/A _7462_/A VGND VGND VPWR VPWR _6576_/B sky130_fd_sc_hd__nand2_1
X_8314_ _8312_/Y _8313_/X _8171_/X _8210_/B VGND VGND VPWR VPWR _8325_/A sky130_fd_sc_hd__o211a_1
X_5526_ _5339_/A _5525_/X _5670_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8245_ _6192_/X _8721_/B _8516_/B _8349_/A VGND VGND VPWR VPWR _8245_/Y sky130_fd_sc_hd__a22oi_1
X_5457_ _5402_/X _5456_/X _5481_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8176_ _8176_/A _8176_/B VGND VGND VPWR VPWR _8179_/A sky130_fd_sc_hd__nor2_1
X_5388_ _9088_/Q VGND VGND VPWR VPWR _5389_/A sky130_fd_sc_hd__clkinv_2
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7127_ _7126_/A _7126_/B _7126_/C VGND VGND VPWR VPWR _7139_/C sky130_fd_sc_hd__a21o_2
X_7058_ _7058_/A _7075_/C VGND VGND VPWR VPWR _7073_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6009_ _6010_/A _6010_/B _6010_/C VGND VGND VPWR VPWR _6018_/B sky130_fd_sc_hd__a21o_1
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4690_ _4701_/A VGND VGND VPWR VPWR _4837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6360_ _7081_/A _6361_/C _7610_/B _6567_/B VGND VGND VPWR VPWR _6362_/A sky130_fd_sc_hd__a22oi_2
X_5311_ _9070_/Q _5337_/B VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__or2_1
X_8030_ _8029_/A _8029_/B _8028_/Y VGND VGND VPWR VPWR _8031_/B sky130_fd_sc_hd__o21ba_1
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6291_ _6292_/B _6378_/A _6292_/A VGND VGND VPWR VPWR _6293_/A sky130_fd_sc_hd__a21o_1
X_5242_ _9068_/Q _5337_/B VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__or2_1
X_5173_ _5173_/A VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 A[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
X_8932_ _8932_/A _8932_/B VGND VGND VPWR VPWR _8935_/A sky130_fd_sc_hd__xor2_1
XFILLER_45_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8863_ _8863_/A _8807_/B VGND VGND VPWR VPWR _8865_/C sky130_fd_sc_hd__or2b_1
X_7814_ _7918_/A _8044_/B VGND VGND VPWR VPWR _7816_/B sky130_fd_sc_hd__and2_1
XFILLER_101_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8794_ _8909_/A _8794_/B VGND VGND VPWR VPWR _8795_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7745_ _7745_/A _7745_/B _7745_/C VGND VGND VPWR VPWR _7746_/B sky130_fd_sc_hd__and3_1
X_4957_ _4957_/A _4957_/B VGND VGND VPWR VPWR _4957_/Y sky130_fd_sc_hd__nor2_1
X_7676_ _7677_/B _7677_/C _7677_/A VGND VGND VPWR VPWR _7796_/B sky130_fd_sc_hd__a21oi_4
X_4888_ _4541_/X _4850_/B _4885_/X _4887_/Y _4889_/A VGND VGND VPWR VPWR _4888_/X
+ sky130_fd_sc_hd__a221o_1
X_6627_ _8190_/C VGND VGND VPWR VPWR _8542_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6558_ _6560_/A _6560_/B _6653_/A _6557_/X VGND VGND VPWR VPWR _6558_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5509_ _5509_/A VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__clkbuf_2
X_6489_ _6489_/A _6432_/B VGND VGND VPWR VPWR _6508_/B sky130_fd_sc_hd__or2b_1
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8228_ _8229_/A _8229_/B _8229_/C VGND VGND VPWR VPWR _8230_/A sky130_fd_sc_hd__a21oi_2
X_8159_ _8159_/A _8159_/B VGND VGND VPWR VPWR _8236_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5860_ _5858_/X _5860_/B VGND VGND VPWR VPWR _5861_/B sky130_fd_sc_hd__and2b_1
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4811_ _4897_/A VGND VGND VPWR VPWR _5785_/S sky130_fd_sc_hd__clkbuf_2
X_5791_ _6240_/A VGND VGND VPWR VPWR _6151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7530_ _7528_/X _7386_/X _7526_/X _7665_/B VGND VGND VPWR VPWR _7668_/A sky130_fd_sc_hd__a211oi_4
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4742_ _9112_/Q VGND VGND VPWR VPWR _4896_/A sky130_fd_sc_hd__clkbuf_2
X_7461_ _7461_/A _7461_/B VGND VGND VPWR VPWR _7473_/A sky130_fd_sc_hd__xnor2_2
X_4673_ _5173_/A VGND VGND VPWR VPWR _5385_/A sky130_fd_sc_hd__clkbuf_2
X_9200_ _9220_/CLK _9200_/D VGND VGND VPWR VPWR _9200_/Q sky130_fd_sc_hd__dfxtp_4
X_6412_ _6411_/A _6411_/B _6411_/C VGND VGND VPWR VPWR _6483_/B sky130_fd_sc_hd__o21a_1
X_7392_ _7192_/B _7392_/B VGND VGND VPWR VPWR _7392_/X sky130_fd_sc_hd__and2b_1
X_9131_ _9223_/CLK _9131_/D VGND VGND VPWR VPWR _9131_/Q sky130_fd_sc_hd__dfxtp_1
X_6343_ _6342_/A _6342_/B _6342_/C VGND VGND VPWR VPWR _6411_/A sky130_fd_sc_hd__o21a_1
XFILLER_88_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6274_ _6759_/C VGND VGND VPWR VPWR _7852_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9062_ _9062_/A _9062_/B VGND VGND VPWR VPWR _9069_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8013_ _8013_/A _7901_/A VGND VGND VPWR VPWR _8013_/X sky130_fd_sc_hd__or2b_1
X_5225_ _5214_/X _5166_/Y _5223_/X _5224_/Y _4556_/A VGND VGND VPWR VPWR _5225_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5156_ _5156_/A VGND VGND VPWR VPWR _5156_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5087_ _4770_/X _5083_/X _5086_/Y _5739_/S VGND VGND VPWR VPWR _5087_/X sky130_fd_sc_hd__o211a_1
X_8915_ _8916_/A _8963_/A _8914_/Y VGND VGND VPWR VPWR _8918_/A sky130_fd_sc_hd__o21a_1
XFILLER_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8846_ _8949_/A _8846_/B VGND VGND VPWR VPWR _8847_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8777_ _8750_/A _8777_/B VGND VGND VPWR VPWR _8819_/A sky130_fd_sc_hd__and2b_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _5990_/B _5989_/B VGND VGND VPWR VPWR _6041_/A sky130_fd_sc_hd__and2b_1
X_7728_ _7938_/B _7728_/B _7728_/C _7728_/D VGND VGND VPWR VPWR _7729_/B sky130_fd_sc_hd__and4_1
XFILLER_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _9198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7659_ _7780_/B _7659_/B VGND VGND VPWR VPWR _7660_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_61 _8438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5010_ _4786_/S _5050_/B _5009_/X VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__a21o_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8700_ _8700_/A _8756_/B VGND VGND VPWR VPWR _8701_/B sky130_fd_sc_hd__nand2_1
X_6961_ _6961_/A _6961_/B VGND VGND VPWR VPWR _6988_/B sky130_fd_sc_hd__or2_2
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6892_ _6892_/A _7022_/B VGND VGND VPWR VPWR _6994_/A sky130_fd_sc_hd__nor2_1
X_5912_ _6660_/A _6825_/B VGND VGND VPWR VPWR _5913_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8631_ _8631_/A _8694_/A _8631_/C VGND VGND VPWR VPWR _8705_/A sky130_fd_sc_hd__or3_2
X_5843_ _6256_/A _6240_/A _5908_/B _5985_/A VGND VGND VPWR VPWR _5844_/B sky130_fd_sc_hd__and4_1
X_8562_ _8562_/A _8631_/A _8562_/C VGND VGND VPWR VPWR _8571_/B sky130_fd_sc_hd__and3_1
X_7513_ _7513_/A _7513_/B VGND VGND VPWR VPWR _7514_/C sky130_fd_sc_hd__xor2_1
X_5774_ _5765_/A _5773_/X _5673_/S VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__o21a_1
X_8493_ _8498_/A _8933_/B _8377_/A _8492_/X VGND VGND VPWR VPWR _8494_/C sky130_fd_sc_hd__a31oi_1
X_4725_ _4721_/X _4693_/Y _4724_/X VGND VGND VPWR VPWR _4725_/Y sky130_fd_sc_hd__a21oi_1
X_7444_ _7445_/A _7445_/B VGND VGND VPWR VPWR _7446_/A sky130_fd_sc_hd__nand2_1
X_4656_ _4656_/A _9107_/Q VGND VGND VPWR VPWR _4676_/B sky130_fd_sc_hd__or2_1
X_7375_ _7518_/A _7518_/B _7518_/C VGND VGND VPWR VPWR _7375_/X sky130_fd_sc_hd__and3_1
X_4587_ _4661_/A VGND VGND VPWR VPWR _4587_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_9114_ _9222_/CLK hold5/X VGND VGND VPWR VPWR _9114_/Q sky130_fd_sc_hd__dfxtp_2
X_6326_ _7770_/A _7453_/A _7457_/A _7647_/A VGND VGND VPWR VPWR _6327_/B sky130_fd_sc_hd__a22oi_2
XFILLER_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9045_ _9045_/A _9045_/B VGND VGND VPWR VPWR _9046_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6257_ _6405_/B _7199_/A _6257_/C _6907_/B VGND VGND VPWR VPWR _6258_/B sky130_fd_sc_hd__and4_1
X_6188_ _9203_/Q VGND VGND VPWR VPWR _7152_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5208_ _5208_/A VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__buf_2
X_5139_ _9074_/Q VGND VGND VPWR VPWR _5430_/A sky130_fd_sc_hd__buf_2
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8829_ _8829_/A _8829_/B VGND VGND VPWR VPWR _8878_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5490_ _5138_/X _5273_/X _5158_/X VGND VGND VPWR VPWR _5490_/Y sky130_fd_sc_hd__a21oi_1
X_7160_ _7160_/A _7160_/B VGND VGND VPWR VPWR _7161_/C sky130_fd_sc_hd__or2_1
XFILLER_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6111_ _7042_/B VGND VGND VPWR VPWR _6361_/C sky130_fd_sc_hd__buf_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _6567_/B _7694_/C _7923_/D _6858_/A VGND VGND VPWR VPWR _7094_/A sky130_fd_sc_hd__a22oi_1
XFILLER_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6040_/Y _6041_/X _5997_/B _5999_/A VGND VGND VPWR VPWR _6044_/C sky130_fd_sc_hd__o211ai_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7993_ _7993_/A _7993_/B VGND VGND VPWR VPWR _8100_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6944_ _6944_/A _6960_/B _6944_/C _7059_/A VGND VGND VPWR VPWR _7059_/B sky130_fd_sc_hd__nor4_2
X_8614_ _8614_/A _8614_/B _8614_/C VGND VGND VPWR VPWR _8615_/B sky130_fd_sc_hd__or3_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6875_ _6875_/A _8844_/A VGND VGND VPWR VPWR _6877_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5826_ _7509_/A _6361_/B _5870_/B _5825_/X VGND VGND VPWR VPWR _5834_/B sky130_fd_sc_hd__a31o_1
XFILLER_22_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8545_ _8677_/A _8782_/A _8545_/C VGND VGND VPWR VPWR _8614_/B sky130_fd_sc_hd__and3_1
X_5757_ _5315_/A _5618_/X _5402_/A _4872_/S VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__o31a_1
X_8476_ _8477_/A _8477_/B VGND VGND VPWR VPWR _8478_/A sky130_fd_sc_hd__nand2_1
X_4708_ _4705_/A _4706_/X _4857_/A VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__mux2_1
X_7427_ _7428_/A _7428_/B VGND VGND VPWR VPWR _7429_/A sky130_fd_sc_hd__nor2_1
X_5688_ _4786_/S _9101_/Q _9102_/Q VGND VGND VPWR VPWR _5688_/Y sky130_fd_sc_hd__a21oi_1
X_4639_ _5227_/A VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7358_ _6151_/A _9184_/Q _7503_/C VGND VGND VPWR VPWR _7358_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ _7040_/A VGND VGND VPWR VPWR _6679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7289_ _7289_/A _7289_/B VGND VGND VPWR VPWR _7552_/B sky130_fd_sc_hd__xor2_2
X_9028_ _9028_/A _9028_/B VGND VGND VPWR VPWR _9029_/C sky130_fd_sc_hd__nor2_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4990_ _4991_/A _4991_/B VGND VGND VPWR VPWR _4992_/A sky130_fd_sc_hd__and2_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6660_ _6660_/A _7822_/B VGND VGND VPWR VPWR _6665_/A sky130_fd_sc_hd__nand2_1
X_6591_ _6591_/A _6591_/B VGND VGND VPWR VPWR _6592_/B sky130_fd_sc_hd__nor2_1
X_5611_ _5368_/X _5119_/A _5609_/X _5610_/Y _5156_/X VGND VGND VPWR VPWR _5611_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8330_ _8331_/A _8331_/B _8329_/Y VGND VGND VPWR VPWR _8510_/A sky130_fd_sc_hd__o21ba_1
X_5542_ _5247_/X _5389_/X _4558_/A VGND VGND VPWR VPWR _5542_/Y sky130_fd_sc_hd__a21oi_1
X_8261_ _8926_/B VGND VGND VPWR VPWR _8978_/B sky130_fd_sc_hd__buf_2
X_5473_ _4721_/X _5420_/X _5471_/X _5472_/Y _5230_/X VGND VGND VPWR VPWR _5473_/X
+ sky130_fd_sc_hd__a221o_1
X_8192_ _8268_/A _8467_/A _8193_/C VGND VGND VPWR VPWR _8194_/A sky130_fd_sc_hd__a21oi_1
X_7212_ _7164_/A _7212_/B _7212_/C VGND VGND VPWR VPWR _7212_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7143_ _7046_/B _7143_/B VGND VGND VPWR VPWR _7143_/X sky130_fd_sc_hd__and2b_1
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ _7061_/A _7061_/B _7073_/X VGND VGND VPWR VPWR _7177_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6025_/A _9163_/Q _7349_/A _7019_/B VGND VGND VPWR VPWR _6029_/A sky130_fd_sc_hd__and4_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7976_ _7976_/A _7976_/B _7976_/C VGND VGND VPWR VPWR _7976_/Y sky130_fd_sc_hd__nand3_2
XFILLER_42_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6927_ _7325_/A _7706_/A _6927_/C _6927_/D VGND VGND VPWR VPWR _6929_/A sky130_fd_sc_hd__and4_1
XFILLER_35_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6858_ _6858_/A _7309_/B VGND VGND VPWR VPWR _6862_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5809_ _7367_/A _7367_/B _6025_/A VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__and3_1
X_8528_ _8538_/A _8792_/B _8792_/D _8530_/A VGND VGND VPWR VPWR _8532_/D sky130_fd_sc_hd__a22o_1
X_6789_ _6894_/A _7346_/B _7347_/B _7006_/B VGND VGND VPWR VPWR _6790_/B sky130_fd_sc_hd__a22oi_1
XFILLER_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8459_ _8568_/A _8898_/B VGND VGND VPWR VPWR _8460_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7830_ _7830_/A _7830_/B _7829_/X VGND VGND VPWR VPWR _7832_/A sky130_fd_sc_hd__or3b_1
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7761_ _7761_/A _7761_/B VGND VGND VPWR VPWR _7861_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4973_ _4770_/X _4936_/Y _4937_/X _5103_/A VGND VGND VPWR VPWR _4973_/X sky130_fd_sc_hd__a31o_1
X_7692_ _6607_/A _7419_/C _7419_/D _6922_/B VGND VGND VPWR VPWR _7696_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6712_ _6712_/A _6834_/A VGND VGND VPWR VPWR _6817_/B sky130_fd_sc_hd__nand2_1
X_6643_ _6643_/A _6643_/B VGND VGND VPWR VPWR _6643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6574_ _6574_/A _6574_/B VGND VGND VPWR VPWR _6576_/A sky130_fd_sc_hd__nor2_1
X_8313_ _8405_/B _8412_/B _8405_/A VGND VGND VPWR VPWR _8313_/X sky130_fd_sc_hd__o21a_1
X_5525_ _5314_/A _5524_/Y _5572_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
X_8244_ _8349_/C VGND VGND VPWR VPWR _8522_/A sky130_fd_sc_hd__clkbuf_2
X_5456_ _5364_/X _5454_/X _5553_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8175_ _8279_/A _8175_/B _8269_/A _8175_/D VGND VGND VPWR VPWR _8176_/B sky130_fd_sc_hd__and4_1
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5387_ _4880_/A _5206_/X _5384_/X _5386_/Y _4545_/A VGND VGND VPWR VPWR _5387_/X
+ sky130_fd_sc_hd__a221o_1
X_7126_ _7126_/A _7126_/B _7126_/C VGND VGND VPWR VPWR _7139_/B sky130_fd_sc_hd__nand3_1
X_7057_ _7057_/A _7172_/A VGND VGND VPWR VPWR _7075_/C sky130_fd_sc_hd__nand2_1
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6008_ _5965_/B _5965_/C _5965_/A VGND VGND VPWR VPWR _6010_/C sky130_fd_sc_hd__o21bai_1
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7959_/A _8084_/A _8190_/B _7959_/D VGND VGND VPWR VPWR _7960_/B sky130_fd_sc_hd__and4_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5310_ _5245_/X _5309_/X _5336_/S VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__mux2_1
X_6290_ _6207_/C _6210_/B _6287_/Y _6288_/X VGND VGND VPWR VPWR _6378_/A sky130_fd_sc_hd__a211o_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5241_ _5117_/X _5240_/X _5336_/S VGND VGND VPWR VPWR _5241_/X sky130_fd_sc_hd__mux2_1
X_5172_ _5172_/A VGND VGND VPWR VPWR _5485_/A sky130_fd_sc_hd__buf_2
Xinput2 A[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_8931_ _8892_/Y _8895_/B _9002_/A _8842_/X VGND VGND VPWR VPWR _8932_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8862_ _8862_/A _8797_/A VGND VGND VPWR VPWR _8865_/A sky130_fd_sc_hd__or2b_1
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8793_ _8793_/A _8793_/B VGND VGND VPWR VPWR _8795_/A sky130_fd_sc_hd__nor2_1
X_7813_ _7813_/A _7813_/B VGND VGND VPWR VPWR _7816_/A sky130_fd_sc_hd__xor2_1
XFILLER_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7744_ _7745_/B _7745_/C _7745_/A VGND VGND VPWR VPWR _7746_/A sky130_fd_sc_hd__a21oi_1
XFILLER_61_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4956_ _5378_/A _4953_/X _4955_/X VGND VGND VPWR VPWR _4956_/X sky130_fd_sc_hd__o21a_1
X_4887_ _5678_/A _4950_/A _4541_/X VGND VGND VPWR VPWR _4887_/Y sky130_fd_sc_hd__a21oi_1
X_7675_ _7675_/A _7795_/C VGND VGND VPWR VPWR _7677_/A sky130_fd_sc_hd__xor2_2
X_6626_ _8050_/C VGND VGND VPWR VPWR _8190_/C sky130_fd_sc_hd__buf_4
X_6557_ _6557_/A _6560_/C VGND VGND VPWR VPWR _6557_/X sky130_fd_sc_hd__and2_1
XFILLER_20_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5508_ _5484_/X _5365_/X _5366_/X _5505_/X _5507_/X VGND VGND VPWR VPWR _9139_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6488_ _6488_/A _6431_/B VGND VGND VPWR VPWR _6508_/A sky130_fd_sc_hd__or2b_1
X_8227_ _8234_/A _8234_/B VGND VGND VPWR VPWR _8229_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5439_ _5138_/X _5212_/X _5158_/X VGND VGND VPWR VPWR _5439_/Y sky130_fd_sc_hd__a21oi_1
X_8158_ _8351_/C _8607_/C VGND VGND VPWR VPWR _8159_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7109_/A _7011_/A VGND VGND VPWR VPWR _7126_/A sky130_fd_sc_hd__or2b_1
XFILLER_101_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8089_ _8089_/A _8089_/B VGND VGND VPWR VPWR _8098_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _4810_/A VGND VGND VPWR VPWR _9154_/D sky130_fd_sc_hd__buf_4
X_5790_ _6235_/A VGND VGND VPWR VPWR _6240_/A sky130_fd_sc_hd__buf_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4741_ _4891_/A _4966_/B _4738_/X _4740_/Y _4535_/A VGND VGND VPWR VPWR _4741_/Y
+ sky130_fd_sc_hd__a221oi_1
X_7460_ _7460_/A _7460_/B VGND VGND VPWR VPWR _7461_/B sky130_fd_sc_hd__nor2_1
X_4672_ _4672_/A VGND VGND VPWR VPWR _5173_/A sky130_fd_sc_hd__buf_2
X_6411_ _6411_/A _6411_/B _6411_/C VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__or3_1
X_9130_ _9222_/CLK _9130_/D VGND VGND VPWR VPWR _9130_/Q sky130_fd_sc_hd__dfxtp_1
X_7391_ _8798_/B VGND VGND VPWR VPWR _8850_/B sky130_fd_sc_hd__buf_4
X_6342_ _6342_/A _6342_/B _6342_/C VGND VGND VPWR VPWR _6344_/A sky130_fd_sc_hd__nor3_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6273_ _7152_/A VGND VGND VPWR VPWR _6759_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_9061_ _5948_/A _5948_/B _9064_/A VGND VGND VPWR VPWR _9062_/B sky130_fd_sc_hd__a21oi_1
X_8012_ _8012_/A _8012_/B VGND VGND VPWR VPWR _8122_/A sky130_fd_sc_hd__xnor2_1
X_5224_ _5158_/A _5482_/A _5135_/A VGND VGND VPWR VPWR _5224_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5155_ _9073_/Q VGND VGND VPWR VPWR _5316_/A sky130_fd_sc_hd__inv_2
XFILLER_96_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5086_ _5105_/B _5086_/B VGND VGND VPWR VPWR _5086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8914_ _8867_/A _8949_/B _8868_/A _8866_/A VGND VGND VPWR VPWR _8914_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_25_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8845_ _8845_/A _8845_/B VGND VGND VPWR VPWR _8847_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8776_ _8776_/A _8776_/B VGND VGND VPWR VPWR _8825_/B sky130_fd_sc_hd__nand2_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5988_ _7361_/C _7093_/B _5910_/X _5987_/Y VGND VGND VPWR VPWR _5989_/B sky130_fd_sc_hd__a31o_1
X_7727_ _7604_/C _7728_/C _7847_/C _7604_/B VGND VGND VPWR VPWR _7729_/A sky130_fd_sc_hd__a22oi_1
X_4939_ _4939_/A _4939_/B VGND VGND VPWR VPWR _4940_/C sky130_fd_sc_hd__or2_2
X_7658_ _7658_/A _7658_/B VGND VGND VPWR VPWR _7659_/B sky130_fd_sc_hd__nor2_1
XANTENNA_40 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _9147_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _7784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6695_/A _6609_/B VGND VGND VPWR VPWR _6611_/C sky130_fd_sc_hd__xnor2_1
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7589_ _7589_/A _7589_/B VGND VGND VPWR VPWR _7592_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6960_ _6960_/A _6960_/B VGND VGND VPWR VPWR _7061_/A sky130_fd_sc_hd__or2_2
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5911_ _5987_/A _5987_/B _5910_/X VGND VGND VPWR VPWR _5913_/A sky130_fd_sc_hd__o21a_1
X_6891_ _6891_/A _6891_/B _6891_/C VGND VGND VPWR VPWR _7022_/B sky130_fd_sc_hd__and3_1
XFILLER_19_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8630_ _8694_/A _8631_/C _8631_/A VGND VGND VPWR VPWR _8632_/A sky130_fd_sc_hd__o21ai_1
X_5842_ _7083_/B _7359_/A _6530_/B _5985_/A VGND VGND VPWR VPWR _5844_/A sky130_fd_sc_hd__a22oi_1
X_8561_ _8631_/A _8562_/C _8562_/A VGND VGND VPWR VPWR _8571_/A sky130_fd_sc_hd__a21oi_2
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _5606_/A _5772_/X _5236_/S VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7512_ _7512_/A _7512_/B VGND VGND VPWR VPWR _7513_/B sky130_fd_sc_hd__xnor2_1
X_4724_ _5734_/S _4723_/X _4698_/X _9104_/Q VGND VGND VPWR VPWR _4724_/X sky130_fd_sc_hd__a31o_1
X_8492_ _8375_/B _8492_/B VGND VGND VPWR VPWR _8492_/X sky130_fd_sc_hd__and2b_1
X_7443_ _7443_/A _7443_/B VGND VGND VPWR VPWR _7445_/B sky130_fd_sc_hd__xnor2_1
X_4655_ _5175_/A VGND VGND VPWR VPWR _4656_/A sky130_fd_sc_hd__clkbuf_2
X_7374_ _7373_/A _7373_/B _7373_/C VGND VGND VPWR VPWR _7518_/C sky130_fd_sc_hd__a21o_2
X_4586_ _4586_/A VGND VGND VPWR VPWR _4661_/A sky130_fd_sc_hd__clkbuf_2
Xinput60 B[5] VGND VGND VPWR VPWR _9198_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_89_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6325_ _6325_/A _6325_/B _7153_/C _7822_/A VGND VGND VPWR VPWR _6327_/A sky130_fd_sc_hd__and4_1
X_9113_ _9199_/CLK hold8/X VGND VGND VPWR VPWR _9113_/Q sky130_fd_sc_hd__dfxtp_4
X_9044_ _9029_/B _8989_/B _9031_/A VGND VGND VPWR VPWR _9045_/B sky130_fd_sc_hd__a21oi_1
XFILLER_88_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6256_ _6256_/A VGND VGND VPWR VPWR _7199_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5207_ _9085_/Q VGND VGND VPWR VPWR _5208_/A sky130_fd_sc_hd__buf_2
X_6187_ _6187_/A _6102_/B VGND VGND VPWR VPWR _6204_/B sky130_fd_sc_hd__or2b_1
XFILLER_96_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5138_ _5156_/A VGND VGND VPWR VPWR _5138_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5069_ _4957_/A _4957_/B _5067_/X _5068_/Y VGND VGND VPWR VPWR _5069_/X sky130_fd_sc_hd__a31o_1
XFILLER_72_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8828_ _8880_/B _8828_/B VGND VGND VPWR VPWR _9104_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8759_ _8759_/A _8759_/B VGND VGND VPWR VPWR _8819_/B sky130_fd_sc_hd__and2_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6110_ _9202_/Q VGND VGND VPWR VPWR _7042_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _9211_/Q VGND VGND VPWR VPWR _7694_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_98_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6041_/A _6041_/B _6041_/C VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__and3_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7992_ _7993_/A _7993_/B VGND VGND VPWR VPWR _7994_/A sky130_fd_sc_hd__or2_1
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6943_ _6944_/A _6960_/B _6944_/C _7059_/A VGND VGND VPWR VPWR _6943_/X sky130_fd_sc_hd__o22a_1
X_6874_ _8595_/C VGND VGND VPWR VPWR _8844_/A sky130_fd_sc_hd__buf_4
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8613_ _8614_/A _8614_/B _8614_/C VGND VGND VPWR VPWR _8672_/B sky130_fd_sc_hd__o21ai_1
XFILLER_62_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5825_ _7006_/A _7506_/B _5940_/A _6031_/A VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__and4_1
X_8544_ _8677_/A _8666_/A _8545_/C VGND VGND VPWR VPWR _8546_/A sky130_fd_sc_hd__a21oi_1
X_5756_ _4676_/B _5755_/X _5282_/S VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__o21a_1
X_8475_ _8392_/A _8392_/B _8474_/X VGND VGND VPWR VPWR _8477_/B sky130_fd_sc_hd__a21oi_1
X_5687_ _5151_/A _5000_/A _5685_/X _5686_/Y _9101_/Q VGND VGND VPWR VPWR _5687_/X
+ sky130_fd_sc_hd__a221o_1
X_4707_ _9095_/Q VGND VGND VPWR VPWR _4857_/A sky130_fd_sc_hd__inv_2
X_7426_ _7562_/A _9214_/Q VGND VGND VPWR VPWR _7428_/B sky130_fd_sc_hd__and2_1
X_4638_ _9102_/Q VGND VGND VPWR VPWR _5227_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7357_ _7357_/A _7357_/B VGND VGND VPWR VPWR _7373_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4569_ _4706_/S VGND VGND VPWR VPWR _4570_/A sky130_fd_sc_hd__buf_2
X_6308_ _7767_/A _7925_/A VGND VGND VPWR VPWR _6321_/A sky130_fd_sc_hd__nand2_2
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7288_ _7405_/A _7288_/B VGND VGND VPWR VPWR _7289_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9027_ _9027_/A _9027_/B VGND VGND VPWR VPWR _9028_/B sky130_fd_sc_hd__and2_1
X_6239_ _7152_/D VGND VGND VPWR VPWR _7455_/A sky130_fd_sc_hd__buf_2
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6590_ _7016_/A _6590_/B _7455_/A _7610_/D VGND VGND VPWR VPWR _6591_/B sky130_fd_sc_hd__and4_1
X_5610_ _5142_/X _5194_/X _5368_/A VGND VGND VPWR VPWR _5610_/Y sky130_fd_sc_hd__a21oi_1
X_5541_ _5160_/X _5205_/A _5539_/X _5540_/Y _5410_/X VGND VGND VPWR VPWR _5541_/X
+ sky130_fd_sc_hd__a221o_1
X_8260_ _8832_/B VGND VGND VPWR VPWR _8926_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_105_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5472_ _4723_/X _5120_/A _4672_/A VGND VGND VPWR VPWR _5472_/Y sky130_fd_sc_hd__a21oi_1
X_7211_ _7321_/A _7321_/B VGND VGND VPWR VPWR _7211_/Y sky130_fd_sc_hd__nor2_1
X_8191_ _8191_/A _8299_/A VGND VGND VPWR VPWR _8193_/C sky130_fd_sc_hd__nor2_1
X_7142_ _7141_/A _7141_/B _7141_/C VGND VGND VPWR VPWR _7218_/A sky130_fd_sc_hd__a21oi_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7073_ _7060_/B _7073_/B VGND VGND VPWR VPWR _7073_/X sky130_fd_sc_hd__and2b_1
XFILLER_100_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6024_ _9200_/Q VGND VGND VPWR VPWR _7019_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7975_ _7975_/A _7975_/B VGND VGND VPWR VPWR _7976_/C sky130_fd_sc_hd__or2_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6926_ _7694_/B _7462_/A VGND VGND VPWR VPWR _6930_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6857_ _9210_/Q VGND VGND VPWR VPWR _7309_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6788_ _9176_/Q VGND VGND VPWR VPWR _7346_/B sky130_fd_sc_hd__clkbuf_2
X_5808_ _9164_/Q VGND VGND VPWR VPWR _6025_/A sky130_fd_sc_hd__clkbuf_2
X_8527_ _8527_/A VGND VGND VPWR VPWR _8700_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5739_ _4545_/A _5738_/X _5739_/S VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8458_ _8563_/B _8458_/B VGND VGND VPWR VPWR _8460_/A sky130_fd_sc_hd__xnor2_1
X_8389_ _8597_/A _8782_/A VGND VGND VPWR VPWR _8390_/B sky130_fd_sc_hd__nand2_1
X_7409_ _7408_/B _7408_/C _7408_/A VGND VGND VPWR VPWR _7548_/B sky130_fd_sc_hd__o21a_1
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7760_ _7761_/A _7761_/B VGND VGND VPWR VPWR _7762_/A sky130_fd_sc_hd__or2_1
X_4972_ _4972_/A VGND VGND VPWR VPWR _4972_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7691_ _7691_/A _7691_/B VGND VGND VPWR VPWR _7784_/B sky130_fd_sc_hd__nor2_1
X_6711_ _6710_/A _6710_/B _6710_/C VGND VGND VPWR VPWR _6834_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6642_ _6643_/A _6643_/B VGND VGND VPWR VPWR _6642_/X sky130_fd_sc_hd__or2_1
X_8312_ _8405_/A _8405_/B _8412_/B VGND VGND VPWR VPWR _8312_/Y sky130_fd_sc_hd__nor3_1
X_6573_ _6922_/B _6927_/C _6927_/D _6754_/B VGND VGND VPWR VPWR _6574_/B sky130_fd_sc_hd__a22oi_1
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5524_ _5450_/X _4966_/A _5523_/X VGND VGND VPWR VPWR _5524_/Y sky130_fd_sc_hd__o21ai_1
X_8243_ _8243_/A _8243_/B VGND VGND VPWR VPWR _8349_/C sky130_fd_sc_hd__and2_1
X_5455_ _5697_/S VGND VGND VPWR VPWR _5553_/S sky130_fd_sc_hd__clkbuf_2
X_8174_ _8371_/A _8595_/C _8595_/D _8279_/A VGND VGND VPWR VPWR _8176_/A sky130_fd_sc_hd__a22oi_1
XFILLER_99_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7125_ _7251_/A _7251_/B VGND VGND VPWR VPWR _7126_/C sky130_fd_sc_hd__xnor2_1
X_5386_ _5385_/X _5278_/X _4656_/A VGND VGND VPWR VPWR _5386_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7056_ _7054_/Y _6939_/X _7052_/X _7053_/Y VGND VGND VPWR VPWR _7172_/A sky130_fd_sc_hd__a211o_1
X_6007_ _6007_/A _6007_/B _6007_/C VGND VGND VPWR VPWR _6010_/B sky130_fd_sc_hd__nand3_1
XFILLER_54_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _8084_/A _8190_/B _8086_/C _8086_/A VGND VGND VPWR VPWR _7960_/A sky130_fd_sc_hd__a22oi_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7889_ _7889_/A _7889_/B VGND VGND VPWR VPWR _7890_/B sky130_fd_sc_hd__nand2_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A _6909_/B VGND VGND VPWR VPWR _6910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5240_ _5120_/X _5239_/X _5282_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
X_5171_ _9079_/Q VGND VGND VPWR VPWR _5172_/A sky130_fd_sc_hd__inv_2
X_8930_ _8930_/A _8979_/B VGND VGND VPWR VPWR _8932_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 A[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
X_8861_ _8861_/A VGND VGND VPWR VPWR _8870_/A sky130_fd_sc_hd__inv_2
XFILLER_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8792_ _8792_/A _8792_/B _8844_/B _8792_/D VGND VGND VPWR VPWR _8793_/B sky130_fd_sc_hd__and4_1
X_7812_ _7918_/A _8039_/A _7696_/D _7694_/X VGND VGND VPWR VPWR _7813_/B sky130_fd_sc_hd__a31o_1
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7743_ _7615_/A _7615_/B _7742_/X VGND VGND VPWR VPWR _7745_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4955_ _5065_/A _4920_/A _4954_/Y VGND VGND VPWR VPWR _4955_/X sky130_fd_sc_hd__a21o_1
X_4886_ _5403_/A VGND VGND VPWR VPWR _5678_/A sky130_fd_sc_hd__clkbuf_2
X_7674_ _7543_/A _7543_/B _7542_/B VGND VGND VPWR VPWR _7795_/C sky130_fd_sc_hd__o21ai_2
X_6625_ _7706_/C VGND VGND VPWR VPWR _8050_/C sky130_fd_sc_hd__clkbuf_2
X_6556_ _6557_/A _6560_/C VGND VGND VPWR VPWR _6653_/A sky130_fd_sc_hd__nor2_1
X_5507_ _5507_/A _5604_/B VGND VGND VPWR VPWR _5507_/X sky130_fd_sc_hd__or2_1
X_8226_ _8226_/A _8233_/B VGND VGND VPWR VPWR _8234_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6487_ _6487_/A _6487_/B VGND VGND VPWR VPWR _6622_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5438_ _4634_/A _5604_/A _5437_/X _4593_/A VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__a211o_1
X_8157_ _8157_/A _8157_/B VGND VGND VPWR VPWR _8159_/A sky130_fd_sc_hd__nor2_1
X_5369_ _5369_/A VGND VGND VPWR VPWR _5634_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8088_ _8290_/A _8519_/A VGND VGND VPWR VPWR _8089_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7108_ _7106_/X _6987_/B _7104_/X _7281_/B VGND VGND VPWR VPWR _7281_/C sky130_fd_sc_hd__a211oi_2
XFILLER_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7039_ _7039_/A _7039_/B VGND VGND VPWR VPWR _7047_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4740_ _4737_/X _4705_/A _4739_/X VGND VGND VPWR VPWR _4740_/Y sky130_fd_sc_hd__a21oi_1
X_4671_ _4721_/A VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7390_ _8044_/B VGND VGND VPWR VPWR _8798_/B sky130_fd_sc_hd__buf_2
X_6410_ _6486_/A _6410_/B VGND VGND VPWR VPWR _6411_/C sky130_fd_sc_hd__xnor2_1
X_6341_ _6341_/A _6341_/B VGND VGND VPWR VPWR _6342_/C sky130_fd_sc_hd__xnor2_2
X_6272_ _9202_/Q VGND VGND VPWR VPWR _7152_/A sky130_fd_sc_hd__clkbuf_2
X_9060_ _9060_/A _9060_/B _9059_/X VGND VGND VPWR VPWR _9070_/D sky130_fd_sc_hd__nor3b_1
X_8011_ _8011_/A _8118_/A VGND VGND VPWR VPWR _8012_/B sky130_fd_sc_hd__xnor2_1
X_5223_ _5215_/X _5370_/A _5220_/X _5221_/Y _5222_/X VGND VGND VPWR VPWR _5223_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5154_ _5154_/A VGND VGND VPWR VPWR _5154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5085_ _4937_/X _5067_/A _5040_/A VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8913_ _8913_/A _8913_/B VGND VGND VPWR VPWR _8963_/A sky130_fd_sc_hd__and2_1
X_8844_ _8844_/A _8844_/B _8844_/C _8844_/D VGND VGND VPWR VPWR _8845_/B sky130_fd_sc_hd__and4_1
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8775_ _8880_/A _8775_/B VGND VGND VPWR VPWR _9103_/D sky130_fd_sc_hd__xnor2_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5987_ _5987_/A _5987_/B VGND VGND VPWR VPWR _5987_/Y sky130_fd_sc_hd__nor2_1
X_7726_ _7726_/A _7637_/A VGND VGND VPWR VPWR _7740_/B sky130_fd_sc_hd__or2b_1
X_4938_ _4939_/A _4939_/B VGND VGND VPWR VPWR _4940_/B sky130_fd_sc_hd__nand2_1
X_7657_ _7657_/A _7657_/B VGND VGND VPWR VPWR _7780_/B sky130_fd_sc_hd__xor2_1
XANTENNA_41 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 _5287_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _5249_/A _4844_/X _4845_/Y _4863_/X _4868_/Y VGND VGND VPWR VPWR _4869_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_52 _9183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _6608_/A _6608_/B VGND VGND VPWR VPWR _6609_/B sky130_fd_sc_hd__xnor2_1
X_7588_ _7588_/A _7714_/B VGND VGND VPWR VPWR _7589_/B sky130_fd_sc_hd__xnor2_1
X_6539_ _6539_/A _6584_/A VGND VGND VPWR VPWR _6585_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8209_ _8209_/A _8209_/B VGND VGND VPWR VPWR _8210_/B sky130_fd_sc_hd__or2_1
X_9189_ _9218_/CLK _9189_/D VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5910_ _7253_/A _6232_/A _7253_/B _6025_/A VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__a22o_1
X_6890_ _6891_/B _6891_/C _6891_/A VGND VGND VPWR VPWR _6892_/A sky130_fd_sc_hd__a21oi_1
X_5841_ _9163_/Q VGND VGND VPWR VPWR _5985_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8560_ _8559_/B _8635_/B _8559_/A VGND VGND VPWR VPWR _8562_/C sky130_fd_sc_hd__o21ai_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5772_ _5557_/A _5771_/X _5714_/S VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__o21a_1
X_7511_ _7369_/A _7368_/A _7368_/B VGND VGND VPWR VPWR _7512_/B sky130_fd_sc_hd__o21ba_1
X_8491_ _8490_/A _8490_/B _8490_/C VGND VGND VPWR VPWR _8501_/B sky130_fd_sc_hd__o21a_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4723_ _5227_/A VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__clkbuf_2
X_7442_ _7312_/A _7312_/B _7441_/X VGND VGND VPWR VPWR _7443_/B sky130_fd_sc_hd__a21oi_1
X_4654_ _4878_/A VGND VGND VPWR VPWR _5175_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7373_ _7373_/A _7373_/B _7373_/C VGND VGND VPWR VPWR _7518_/B sky130_fd_sc_hd__nand3_1
Xinput50 B[25] VGND VGND VPWR VPWR _9218_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 B[6] VGND VGND VPWR VPWR _9199_/D sky130_fd_sc_hd__clkbuf_1
X_4585_ _4585_/A VGND VGND VPWR VPWR _4586_/A sky130_fd_sc_hd__clkbuf_2
X_6324_ _9171_/Q VGND VGND VPWR VPWR _7153_/C sky130_fd_sc_hd__clkbuf_2
X_9112_ _9218_/CLK _9112_/D VGND VGND VPWR VPWR _9112_/Q sky130_fd_sc_hd__dfxtp_2
X_9043_ _8989_/B _9031_/A _9028_/B VGND VGND VPWR VPWR _9045_/A sky130_fd_sc_hd__a21o_1
X_6255_ _6974_/B VGND VGND VPWR VPWR _6405_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5206_ _5206_/A VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__buf_2
XFILLER_88_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6186_ _6186_/A _6101_/B VGND VGND VPWR VPWR _6204_/A sky130_fd_sc_hd__or2b_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5137_ _9076_/Q VGND VGND VPWR VPWR _5482_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5068_ _4957_/A _5046_/B _5074_/B VGND VGND VPWR VPWR _5068_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8827_ _8768_/X _8775_/B _8769_/A VGND VGND VPWR VPWR _8828_/B sky130_fd_sc_hd__a21o_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8758_ _8759_/A _8759_/B VGND VGND VPWR VPWR _8760_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7709_ _7819_/C _7709_/B VGND VGND VPWR VPWR _7818_/B sky130_fd_sc_hd__xnor2_1
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8689_ _8687_/Y _8753_/A _8620_/B _8624_/C VGND VGND VPWR VPWR _8691_/C sky130_fd_sc_hd__o211a_1
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6041_/B _6041_/C _6041_/A VGND VGND VPWR VPWR _6040_/Y sky130_fd_sc_hd__a21oi_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7991_ _7991_/A _8078_/B VGND VGND VPWR VPWR _7993_/B sky130_fd_sc_hd__nor2_1
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6942_ _6940_/D _6940_/Y _6938_/Y _6939_/X VGND VGND VPWR VPWR _7059_/A sky130_fd_sc_hd__o211a_1
X_6873_ _8269_/A VGND VGND VPWR VPWR _8595_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8612_ _8661_/A _8612_/B VGND VGND VPWR VPWR _8614_/C sky130_fd_sc_hd__xnor2_1
X_5824_ _7367_/B VGND VGND VPWR VPWR _7506_/B sky130_fd_sc_hd__buf_2
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8543_ _8543_/A _8614_/A VGND VGND VPWR VPWR _8545_/C sky130_fd_sc_hd__nor2_1
X_5755_ _5509_/X _5583_/X _5750_/X _5754_/X _5676_/A VGND VGND VPWR VPWR _5755_/X
+ sky130_fd_sc_hd__o311a_1
X_8474_ _8391_/A _8474_/B VGND VGND VPWR VPWR _8474_/X sky130_fd_sc_hd__and2b_1
X_5686_ _4571_/A _5002_/A _9100_/Q VGND VGND VPWR VPWR _5686_/Y sky130_fd_sc_hd__a21oi_1
X_4706_ _4759_/A _4705_/Y _4706_/S VGND VGND VPWR VPWR _4706_/X sky130_fd_sc_hd__mux2_1
X_7425_ _7425_/A _7425_/B VGND VGND VPWR VPWR _7428_/A sky130_fd_sc_hd__xor2_1
X_4637_ _4637_/A VGND VGND VPWR VPWR _5534_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7356_ _7356_/A _7263_/A VGND VGND VPWR VPWR _7373_/A sky130_fd_sc_hd__or2b_1
X_4568_ _4568_/A VGND VGND VPWR VPWR _4706_/S sky130_fd_sc_hd__buf_2
X_6307_ _7435_/A VGND VGND VPWR VPWR _7925_/A sky130_fd_sc_hd__clkbuf_2
X_7287_ _7287_/A _7287_/B _7287_/C VGND VGND VPWR VPWR _7288_/B sky130_fd_sc_hd__or3_1
XFILLER_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9026_ _9027_/A _9027_/B VGND VGND VPWR VPWR _9028_/A sky130_fd_sc_hd__nor2_1
X_6238_ _9173_/Q VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A VGND VGND VPWR VPWR _7083_/A sky130_fd_sc_hd__clkbuf_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5540_ _5138_/X _5656_/A _5158_/X VGND VGND VPWR VPWR _5540_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5471_ _5213_/X _5194_/X _5469_/X _5470_/Y _5227_/X VGND VGND VPWR VPWR _5471_/X
+ sky130_fd_sc_hd__a221o_1
X_7210_ _7321_/A _7321_/B VGND VGND VPWR VPWR _7210_/X sky130_fd_sc_hd__and2_1
X_8190_ _8190_/A _8190_/B _8190_/C _8720_/A VGND VGND VPWR VPWR _8299_/A sky130_fd_sc_hd__and4_1
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7141_ _7141_/A _7141_/B _7141_/C VGND VGND VPWR VPWR _7166_/B sky130_fd_sc_hd__and3_2
XFILLER_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7072_ _7072_/A _7072_/B VGND VGND VPWR VPWR _7182_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6023_ _6825_/A _6660_/A _5971_/B _5969_/X VGND VGND VPWR VPWR _6107_/A sky130_fd_sc_hd__a31o_1
XFILLER_100_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7974_ _7974_/A _7974_/B VGND VGND VPWR VPWR _7975_/B sky130_fd_sc_hd__and2_1
XFILLER_66_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6925_ _6925_/A VGND VGND VPWR VPWR _7694_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6856_ _6757_/A _6756_/B _6756_/A VGND VGND VPWR VPWR _6982_/A sky130_fd_sc_hd__o21ba_1
X_6787_ _7259_/A _7259_/B _7131_/D _7347_/B VGND VGND VPWR VPWR _6790_/A sky130_fd_sc_hd__and4_1
X_5807_ _6667_/A VGND VGND VPWR VPWR _7367_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8526_ _8624_/A _8526_/B VGND VGND VPWR VPWR _8559_/A sky130_fd_sc_hd__or2_1
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5738_ _5177_/A _5737_/X _5738_/S VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__mux2_1
X_8457_ _8370_/A _8373_/B _8370_/B VGND VGND VPWR VPWR _8458_/B sky130_fd_sc_hd__o21ba_1
X_5669_ _4600_/A _5668_/X _5692_/S VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__mux2_1
X_8388_ _8530_/A VGND VGND VPWR VPWR _8597_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7408_ _7408_/A _7408_/B _7408_/C VGND VGND VPWR VPWR _7410_/A sky130_fd_sc_hd__nor3_1
XFILLER_89_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7339_ _7339_/A _7339_/B VGND VGND VPWR VPWR _7340_/C sky130_fd_sc_hd__or2_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9009_ _9009_/A _9009_/B _9009_/C VGND VGND VPWR VPWR _9032_/A sky130_fd_sc_hd__and3_1
XFILLER_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4971_ _5670_/S _4971_/B VGND VGND VPWR VPWR _4972_/A sky130_fd_sc_hd__nor2_1
X_7690_ _7690_/A _7690_/B VGND VGND VPWR VPWR _7799_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6710_ _6710_/A _6710_/B _6710_/C VGND VGND VPWR VPWR _6712_/A sky130_fd_sc_hd__nand3_1
X_6641_ _6641_/A _6641_/B VGND VGND VPWR VPWR _6656_/A sky130_fd_sc_hd__nor2_2
X_8311_ _8199_/B _8202_/B _8308_/X _8412_/A VGND VGND VPWR VPWR _8412_/B sky130_fd_sc_hd__a211oi_4
X_6572_ _7199_/A _6572_/B _7042_/B _6572_/D VGND VGND VPWR VPWR _6574_/A sky130_fd_sc_hd__and4_1
X_5523_ _5424_/X _4721_/X _5521_/X _5522_/Y _5230_/X VGND VGND VPWR VPWR _5523_/X
+ sky130_fd_sc_hd__a221o_1
X_8242_ _8242_/A _8242_/B VGND VGND VPWR VPWR _8252_/A sky130_fd_sc_hd__xnor2_1
X_5454_ _5339_/X _5452_/X _5552_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8173_ _8175_/B VGND VGND VPWR VPWR _8371_/A sky130_fd_sc_hd__clkbuf_2
X_5385_ _5385_/A VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7124_ _7124_/A _7250_/A VGND VGND VPWR VPWR _7251_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7055_ _7052_/X _7053_/Y _7054_/Y _6939_/X VGND VGND VPWR VPWR _7057_/A sky130_fd_sc_hd__o211ai_1
XFILLER_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6006_ _6007_/B _6007_/C _6007_/A VGND VGND VPWR VPWR _6010_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7957_ _7957_/A _7878_/A VGND VGND VPWR VPWR _7976_/B sky130_fd_sc_hd__or2b_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7888_ _7888_/A _7887_/A VGND VGND VPWR VPWR _7889_/B sky130_fd_sc_hd__or2b_1
X_6908_ _6908_/A _6908_/B VGND VGND VPWR VPWR _6909_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6839_ _6945_/A _6945_/B _6945_/C VGND VGND VPWR VPWR _6839_/X sky130_fd_sc_hd__and3_1
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8509_ _8580_/A _8580_/B VGND VGND VPWR VPWR _8512_/A sky130_fd_sc_hd__xnor2_2
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5170_ _5414_/A VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 A[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_8860_ _8908_/A _8860_/B VGND VGND VPWR VPWR _8861_/A sky130_fd_sc_hd__and2_1
X_8791_ _8844_/A _8844_/B _8844_/C _8949_/A VGND VGND VPWR VPWR _8793_/A sky130_fd_sc_hd__a22oi_1
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7811_ _7811_/A _7811_/B VGND VGND VPWR VPWR _7813_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7742_ _7614_/B _7742_/B VGND VGND VPWR VPWR _7742_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4954_ _5065_/A _4920_/A _4556_/A VGND VGND VPWR VPWR _4954_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7673_ _7795_/A _7795_/B VGND VGND VPWR VPWR _7675_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4885_ _5714_/S _4881_/X _4882_/Y _4884_/X VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6624_ _9208_/Q VGND VGND VPWR VPWR _7706_/C sky130_fd_sc_hd__clkbuf_2
X_6555_ _6655_/A _6655_/B VGND VGND VPWR VPWR _6560_/C sky130_fd_sc_hd__xnor2_1
X_5506_ _5506_/A VGND VGND VPWR VPWR _5604_/B sky130_fd_sc_hd__clkbuf_1
X_8225_ _8114_/A _8114_/B _8117_/B VGND VGND VPWR VPWR _8233_/B sky130_fd_sc_hd__o21bai_2
X_6486_ _6486_/A _6410_/B VGND VGND VPWR VPWR _6487_/B sky130_fd_sc_hd__or2b_1
X_5437_ _5618_/A _5131_/A _5435_/X _5436_/X _4566_/A VGND VGND VPWR VPWR _5437_/X
+ sky130_fd_sc_hd__o221a_1
X_8156_ _8156_/A _8156_/B _8156_/C _8721_/B VGND VGND VPWR VPWR _8157_/B sky130_fd_sc_hd__and4_1
X_5368_ _5368_/A VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__clkbuf_2
X_8087_ _8087_/A _8087_/B VGND VGND VPWR VPWR _8089_/A sky130_fd_sc_hd__nor2_1
X_5299_ _5385_/A _5184_/X _5175_/A VGND VGND VPWR VPWR _5299_/Y sky130_fd_sc_hd__a21oi_1
X_7107_ _7104_/X _7281_/B _7106_/X _6987_/B VGND VGND VPWR VPWR _7170_/A sky130_fd_sc_hd__o211a_1
XFILLER_101_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7038_ _7038_/A _7038_/B VGND VGND VPWR VPWR _7039_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8989_ _8989_/A _8989_/B VGND VGND VPWR VPWR _8990_/B sky130_fd_sc_hd__nand2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4670_ _5393_/A VGND VGND VPWR VPWR _5200_/A sky130_fd_sc_hd__buf_2
X_6340_ _6340_/A _6340_/B VGND VGND VPWR VPWR _6341_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6271_ _7096_/A _7608_/A VGND VGND VPWR VPWR _6280_/A sky130_fd_sc_hd__nand2_1
X_8010_ _7898_/A _7898_/B _8009_/X VGND VGND VPWR VPWR _8118_/A sky130_fd_sc_hd__a21oi_2
X_5222_ _5222_/A VGND VGND VPWR VPWR _5222_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5153_ _5142_/X _5362_/A _5148_/X _5152_/Y _5368_/A VGND VGND VPWR VPWR _5153_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5084_ _4937_/X _5067_/X _5671_/S VGND VGND VPWR VPWR _5105_/B sky130_fd_sc_hd__a21oi_1
X_8912_ _8913_/A _8913_/B VGND VGND VPWR VPWR _8916_/A sky130_fd_sc_hd__nor2_1
X_8843_ _8989_/A _8450_/D _8842_/X VGND VGND VPWR VPWR _8845_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8774_ _8652_/B _8772_/X _8773_/X _8772_/B VGND VGND VPWR VPWR _8775_/B sky130_fd_sc_hd__a22oi_4
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5986_ _5986_/A _6108_/A VGND VGND VPWR VPWR _5990_/B sky130_fd_sc_hd__or2_1
X_7725_ _7725_/A _7801_/B VGND VGND VPWR VPWR _7783_/A sky130_fd_sc_hd__nor2_1
X_4937_ _4937_/A _4937_/B VGND VGND VPWR VPWR _4937_/X sky130_fd_sc_hd__or2_2
X_7656_ _7776_/B _7656_/B VGND VGND VPWR VPWR _7657_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_20 _9136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4862_/X _4882_/B _5156_/A VGND VGND VPWR VPWR _4868_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_53 _9201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6607_/A _6607_/B VGND VGND VPWR VPWR _6608_/B sky130_fd_sc_hd__nand2_1
XANTENNA_42 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7587_ _7587_/A _7712_/B VGND VGND VPWR VPWR _7714_/B sky130_fd_sc_hd__nor2_1
X_4799_ _4799_/A _4836_/A VGND VGND VPWR VPWR _4799_/Y sky130_fd_sc_hd__nand2_1
X_6538_ _6452_/A _6451_/B _6451_/A VGND VGND VPWR VPWR _6584_/A sky130_fd_sc_hd__o21ba_1
X_6469_ _6469_/A _6469_/B VGND VGND VPWR VPWR _6470_/B sky130_fd_sc_hd__nor2_1
X_9188_ _9208_/CLK _9188_/D VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
X_8208_ _8209_/A _8209_/B VGND VGND VPWR VPWR _8210_/A sky130_fd_sc_hd__nand2_1
X_8139_ _8139_/A _8481_/A VGND VGND VPWR VPWR _8144_/A sky130_fd_sc_hd__and2_1
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5840_ _7253_/B VGND VGND VPWR VPWR _6530_/B sky130_fd_sc_hd__buf_2
XFILLER_61_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5771_ _4560_/A _5770_/X _5712_/S VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7510_ _7645_/C _7510_/B VGND VGND VPWR VPWR _7512_/A sky130_fd_sc_hd__xor2_1
X_8490_ _8490_/A _8490_/B _8490_/C VGND VGND VPWR VPWR _8501_/A sky130_fd_sc_hd__nor3_1
X_4722_ _9103_/Q VGND VGND VPWR VPWR _5734_/S sky130_fd_sc_hd__clkinv_2
X_7441_ _7311_/A _7441_/B VGND VGND VPWR VPWR _7441_/X sky130_fd_sc_hd__and2b_1
Xinput40 B[16] VGND VGND VPWR VPWR _9209_/D sky130_fd_sc_hd__clkbuf_1
X_4653_ _9104_/Q VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__clkbuf_2
X_7372_ _7496_/A _7496_/B VGND VGND VPWR VPWR _7373_/C sky130_fd_sc_hd__xnor2_1
Xinput51 B[26] VGND VGND VPWR VPWR _9219_/D sky130_fd_sc_hd__clkbuf_1
Xinput62 B[7] VGND VGND VPWR VPWR _9200_/D sky130_fd_sc_hd__clkbuf_1
X_4584_ _4584_/A VGND VGND VPWR VPWR _4585_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6323_ _6593_/A _7938_/A VGND VGND VPWR VPWR _6328_/A sky130_fd_sc_hd__nand2_2
X_9111_ _9218_/CLK _9111_/D VGND VGND VPWR VPWR _9111_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9042_ _9032_/A _9032_/B _9041_/Y VGND VGND VPWR VPWR _9046_/A sky130_fd_sc_hd__a21oi_2
X_6254_ _6754_/B _6907_/A _7986_/A _7419_/A VGND VGND VPWR VPWR _6258_/A sky130_fd_sc_hd__a22oi_2
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5205_ _5205_/A VGND VGND VPWR VPWR _5206_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6185_ _6104_/C _6104_/Y _6182_/Y _6183_/X VGND VGND VPWR VPWR _6207_/C sky130_fd_sc_hd__a211o_1
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5136_ _5410_/A VGND VGND VPWR VPWR _5136_/X sky130_fd_sc_hd__clkbuf_2
X_5067_ _5067_/A _5067_/B VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__and2_1
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8826_ _8826_/A _8825_/Y VGND VGND VPWR VPWR _8880_/B sky130_fd_sc_hd__or2b_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8757_ _8757_/A _8757_/B VGND VGND VPWR VPWR _8759_/B sky130_fd_sc_hd__xnor2_1
X_5969_ _9165_/Q _6235_/A _6885_/A _9169_/Q VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__and4_1
X_7708_ _7808_/B _7824_/B VGND VGND VPWR VPWR _7709_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8688_ _8688_/A _8688_/B _8688_/C VGND VGND VPWR VPWR _8753_/A sky130_fd_sc_hd__and3_1
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7639_ _7880_/A _8607_/D _7767_/C VGND VGND VPWR VPWR _7644_/A sky130_fd_sc_hd__a21oi_1
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7990_ _7990_/A _7990_/B _7990_/C VGND VGND VPWR VPWR _8078_/B sky130_fd_sc_hd__and3_1
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6941_ _6938_/Y _6939_/X _6940_/D _6940_/Y VGND VGND VPWR VPWR _6944_/C sky130_fd_sc_hd__a211oi_2
X_6872_ _7923_/C VGND VGND VPWR VPWR _8269_/A sky130_fd_sc_hd__clkbuf_2
X_8611_ _8661_/B _8662_/B VGND VGND VPWR VPWR _8612_/B sky130_fd_sc_hd__nor2_1
X_5823_ _7367_/A VGND VGND VPWR VPWR _7006_/A sky130_fd_sc_hd__buf_2
XFILLER_62_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8542_ _8542_/A _8542_/B _8542_/C _8607_/C VGND VGND VPWR VPWR _8614_/A sky130_fd_sc_hd__and4_1
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5754_ _5754_/A _5754_/B _5754_/C VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__or3_1
X_8473_ _8473_/A _8473_/B VGND VGND VPWR VPWR _8477_/A sky130_fd_sc_hd__xnor2_1
X_5685_ _5313_/A _4789_/A _5683_/X _5684_/Y _5002_/A VGND VGND VPWR VPWR _5685_/X
+ sky130_fd_sc_hd__a221o_1
X_4705_ _4705_/A _4705_/B VGND VGND VPWR VPWR _4705_/Y sky130_fd_sc_hd__xnor2_1
X_7424_ _7562_/A _7810_/B _7295_/D _7293_/X VGND VGND VPWR VPWR _7425_/B sky130_fd_sc_hd__a31o_1
X_4636_ _4636_/A VGND VGND VPWR VPWR _5484_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7355_ _7452_/A _7355_/B VGND VGND VPWR VPWR _7518_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6306_ _7307_/B VGND VGND VPWR VPWR _7435_/A sky130_fd_sc_hd__clkbuf_2
X_4567_ _9094_/Q VGND VGND VPWR VPWR _4568_/A sky130_fd_sc_hd__inv_2
X_7286_ _7287_/A _7287_/B _7287_/C VGND VGND VPWR VPWR _7405_/A sky130_fd_sc_hd__o21ai_2
XFILLER_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9025_ _9025_/A _9025_/B VGND VGND VPWR VPWR _9027_/B sky130_fd_sc_hd__and2_1
X_6237_ _6998_/A _6998_/B _6702_/B _7330_/A VGND VGND VPWR VPWR _6342_/A sky130_fd_sc_hd__and4_2
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6081_/A _6085_/B _6081_/B VGND VGND VPWR VPWR _6267_/A sky130_fd_sc_hd__o21ba_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A VGND VGND VPWR VPWR _5120_/A sky130_fd_sc_hd__buf_2
X_6099_ _6359_/A _7988_/A VGND VGND VPWR VPWR _6100_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8809_ _8809_/A _8809_/B VGND VGND VPWR VPWR _8872_/A sky130_fd_sc_hd__or2_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5470_ _4717_/S _5122_/A _4605_/A VGND VGND VPWR VPWR _5470_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7140_ _7140_/A _7140_/B VGND VGND VPWR VPWR _7141_/C sky130_fd_sc_hd__nand2_1
XFILLER_98_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7071_ _7071_/A _7071_/B _7071_/C VGND VGND VPWR VPWR _7406_/A sky130_fd_sc_hd__nand3_1
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6022_/A VGND VGND VPWR VPWR _6825_/A sky130_fd_sc_hd__clkbuf_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7973_ _7974_/A _7974_/B VGND VGND VPWR VPWR _7975_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6924_ _6924_/A _6924_/B VGND VGND VPWR VPWR _6933_/A sky130_fd_sc_hd__xnor2_2
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _6968_/B _8052_/B _6829_/A _6825_/X VGND VGND VPWR VPWR _6864_/A sky130_fd_sc_hd__a31o_1
X_6786_ _9177_/Q VGND VGND VPWR VPWR _7347_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5806_ _9195_/Q VGND VGND VPWR VPWR _6667_/A sky130_fd_sc_hd__clkbuf_2
X_8525_ _8525_/A _8525_/B _8525_/C VGND VGND VPWR VPWR _8526_/B sky130_fd_sc_hd__and3_1
X_5737_ _5129_/A _5736_/X _5737_/S VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__mux2_1
X_8456_ _8456_/A _8456_/B VGND VGND VPWR VPWR _8563_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7407_ _7289_/A _7182_/Y _7289_/B VGND VGND VPWR VPWR _7408_/C sky130_fd_sc_hd__a21oi_2
X_5668_ _5460_/A _5667_/X _5691_/S VGND VGND VPWR VPWR _5668_/X sky130_fd_sc_hd__mux2_1
X_8387_ _8387_/A _8387_/B VGND VGND VPWR VPWR _8390_/A sky130_fd_sc_hd__nor2_1
X_4619_ _5739_/S VGND VGND VPWR VPWR _5695_/S sky130_fd_sc_hd__buf_2
X_5599_ _5749_/A _5598_/X _5671_/S VGND VGND VPWR VPWR _5599_/X sky130_fd_sc_hd__mux2_1
X_7338_ _7338_/A _7338_/B VGND VGND VPWR VPWR _7339_/B sky130_fd_sc_hd__and2_1
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7269_ _7267_/X _7268_/Y _7139_/C _7140_/B VGND VGND VPWR VPWR _7271_/C sky130_fd_sc_hd__o211ai_4
X_9008_ _9008_/A _9008_/B VGND VGND VPWR VPWR _9009_/C sky130_fd_sc_hd__xor2_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4970_ _5737_/S VGND VGND VPWR VPWR _5670_/S sky130_fd_sc_hd__buf_2
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6640_ _6640_/A _6640_/B _6640_/C VGND VGND VPWR VPWR _6641_/B sky130_fd_sc_hd__and3_1
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6571_ _6571_/A _6571_/B VGND VGND VPWR VPWR _6579_/A sky130_fd_sc_hd__xnor2_2
X_8310_ _8308_/X _8412_/A _8199_/B _8202_/B VGND VGND VPWR VPWR _8405_/B sky130_fd_sc_hd__o211a_1
X_5522_ _5200_/A _4723_/X _4672_/A VGND VGND VPWR VPWR _5522_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8241_ _8584_/A _8677_/A VGND VGND VPWR VPWR _8242_/B sky130_fd_sc_hd__nand2_1
X_5453_ _5696_/S VGND VGND VPWR VPWR _5552_/S sky130_fd_sc_hd__clkbuf_2
X_8172_ _8172_/A _8171_/X VGND VGND VPWR VPWR _8209_/A sky130_fd_sc_hd__or2b_1
X_5384_ _5266_/X _5208_/X _5381_/X _5383_/Y _4550_/A VGND VGND VPWR VPWR _5384_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7123_ _7009_/A _7008_/B _7008_/A VGND VGND VPWR VPWR _7250_/A sky130_fd_sc_hd__o21ba_1
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7054_ _7054_/A VGND VGND VPWR VPWR _7054_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6005_ _9194_/Q _9169_/Q VGND VGND VPWR VPWR _6007_/A sky130_fd_sc_hd__and2_1
XFILLER_94_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _7956_/A _8029_/B VGND VGND VPWR VPWR _8007_/A sky130_fd_sc_hd__or2_1
XFILLER_70_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7887_ _7887_/A _7888_/A VGND VGND VPWR VPWR _7889_/A sky130_fd_sc_hd__or2b_1
X_6907_ _6907_/A _6907_/B _7455_/A _7129_/B VGND VGND VPWR VPWR _6908_/B sky130_fd_sc_hd__and4_1
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ _6945_/B _6945_/C _6945_/A VGND VGND VPWR VPWR _6838_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8508_ _8422_/A _8422_/B _8424_/X VGND VGND VPWR VPWR _8580_/B sky130_fd_sc_hd__a21oi_2
X_6769_ _6708_/B _6769_/B VGND VGND VPWR VPWR _6769_/X sky130_fd_sc_hd__and2b_1
XFILLER_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8439_ _8439_/A _8439_/B VGND VGND VPWR VPWR _8442_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 A[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7810_ _7808_/X _7810_/B _7810_/C _7810_/D VGND VGND VPWR VPWR _7811_/B sky130_fd_sc_hd__and4b_1
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8790_ _8790_/A _8790_/B VGND VGND VPWR VPWR _8803_/A sky130_fd_sc_hd__xnor2_1
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7741_ _7740_/A _7740_/B _7740_/C VGND VGND VPWR VPWR _7745_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4953_ _4925_/Y _4926_/X _4952_/X _4598_/A VGND VGND VPWR VPWR _4953_/X sky130_fd_sc_hd__o22a_1
X_7672_ _7672_/A _7672_/B VGND VGND VPWR VPWR _7795_/B sky130_fd_sc_hd__nand2_1
X_4884_ _5632_/A _4844_/X _4845_/Y _4883_/X VGND VGND VPWR VPWR _4884_/X sky130_fd_sc_hd__a31o_1
X_6623_ _7194_/A VGND VGND VPWR VPWR _7389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6554_ _6470_/A _6470_/B _6469_/B VGND VGND VPWR VPWR _6655_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5505_ _5461_/X _5503_/X _5603_/S VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__mux2_1
X_6485_ _6485_/A _6409_/A VGND VGND VPWR VPWR _6487_/A sky130_fd_sc_hd__or2b_1
X_8224_ _8224_/A _8224_/B VGND VGND VPWR VPWR _8226_/A sky130_fd_sc_hd__or2_1
X_5436_ _5149_/A _5555_/A _4586_/A VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8155_ _6192_/X _8156_/C _8154_/X VGND VGND VPWR VPWR _8157_/A sky130_fd_sc_hd__a21oi_1
X_5367_ _5367_/A VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8086_ _8086_/A _8516_/A _8086_/C _8150_/C VGND VGND VPWR VPWR _8087_/B sky130_fd_sc_hd__and4_1
XFILLER_87_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5298_ _5414_/A _5630_/A _5296_/X _5297_/Y _5129_/A VGND VGND VPWR VPWR _5298_/X
+ sky130_fd_sc_hd__a221o_1
X_7106_ _7106_/A _6984_/B VGND VGND VPWR VPWR _7106_/X sky130_fd_sc_hd__or2b_1
XFILLER_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7037_ _7037_/A _7148_/A _7222_/C _7222_/D VGND VGND VPWR VPWR _7038_/B sky130_fd_sc_hd__and4_1
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8988_ _9015_/B _8988_/B VGND VGND VPWR VPWR _8990_/A sky130_fd_sc_hd__xnor2_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7939_/A _8056_/A VGND VGND VPWR VPWR _8047_/C sky130_fd_sc_hd__nor2_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6270_ _7153_/D VGND VGND VPWR VPWR _7608_/A sky130_fd_sc_hd__buf_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5221_ _5154_/A _9074_/Q _4591_/A VGND VGND VPWR VPWR _5221_/Y sky130_fd_sc_hd__a21oi_1
X_5152_ _5149_/X _5150_/Y _5151_/X VGND VGND VPWR VPWR _5152_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5083_ _5046_/Y _5047_/X _5082_/X _4799_/A VGND VGND VPWR VPWR _5083_/X sky130_fd_sc_hd__o2bb2a_1
X_8911_ _8923_/A _8957_/B VGND VGND VPWR VPWR _8913_/B sky130_fd_sc_hd__xnor2_1
X_8842_ _8842_/A _8842_/B VGND VGND VPWR VPWR _8842_/X sky130_fd_sc_hd__and2_1
XFILLER_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8773_ _8773_/A _8773_/B VGND VGND VPWR VPWR _8773_/X sky130_fd_sc_hd__or2_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7724_ _7724_/A _7724_/B _7724_/C VGND VGND VPWR VPWR _7801_/B sky130_fd_sc_hd__and3_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5985_ _5985_/A _9162_/Q _6172_/A _5985_/D VGND VGND VPWR VPWR _6108_/A sky130_fd_sc_hd__and4_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4936_ _4937_/A _4937_/B VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_21 _9136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _9151_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7655_ _7512_/A _7512_/B _7513_/B _7513_/A VGND VGND VPWR VPWR _7656_/B sky130_fd_sc_hd__o22a_1
XANTENNA_32 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _5080_/A _4915_/A VGND VGND VPWR VPWR _4882_/B sky130_fd_sc_hd__or2_2
X_7586_ _7925_/A _7940_/B _7586_/C VGND VGND VPWR VPWR _7712_/B sky130_fd_sc_hd__and3_1
XANTENNA_54 _9212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6606_/A _6606_/B VGND VGND VPWR VPWR _6608_/A sky130_fd_sc_hd__nor2_1
XANTENNA_43 _9195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _6537_/A _6537_/B VGND VGND VPWR VPWR _6539_/A sky130_fd_sc_hd__xnor2_1
X_4798_ _4787_/B _4797_/X _4834_/A VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6468_ _6372_/C _6466_/Y _6551_/B _6465_/X VGND VGND VPWR VPWR _6469_/B sky130_fd_sc_hd__o211a_1
X_9187_ _9210_/CLK _9187_/D VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
X_8207_ _8207_/A _8318_/B VGND VGND VPWR VPWR _8209_/B sky130_fd_sc_hd__or2_1
X_5419_ _9089_/Q VGND VGND VPWR VPWR _5420_/A sky130_fd_sc_hd__inv_2
X_6399_ _6399_/A _6483_/A VGND VGND VPWR VPWR _6486_/A sky130_fd_sc_hd__or2_1
X_8138_ _8257_/C _8138_/B VGND VGND VPWR VPWR _8481_/A sky130_fd_sc_hd__or2_1
XFILLER_101_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8069_ _8069_/A _8720_/B VGND VGND VPWR VPWR _8071_/C sky130_fd_sc_hd__and2_1
XFILLER_75_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A VGND VGND VPWR VPWR _9090_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5770_ _5460_/A _5769_/X _4875_/S VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__o21a_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A VGND VGND VPWR VPWR _4721_/X sky130_fd_sc_hd__clkbuf_2
X_7440_ _7440_/A _7440_/B VGND VGND VPWR VPWR _7443_/A sky130_fd_sc_hd__xnor2_1
X_4652_ _5339_/A _5432_/A _5103_/A _9111_/Q VGND VGND VPWR VPWR _4676_/A sky130_fd_sc_hd__or4_1
Xinput30 A[7] VGND VGND VPWR VPWR _9169_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 B[17] VGND VGND VPWR VPWR _9210_/D sky130_fd_sc_hd__clkbuf_1
Xinput63 B[8] VGND VGND VPWR VPWR _9201_/D sky130_fd_sc_hd__clkbuf_1
X_7371_ _7495_/B _7371_/B VGND VGND VPWR VPWR _7496_/B sky130_fd_sc_hd__xnor2_1
X_9110_ _9218_/CLK _9110_/D VGND VGND VPWR VPWR _9110_/Q sky130_fd_sc_hd__dfxtp_1
Xinput52 B[27] VGND VGND VPWR VPWR _9220_/D sky130_fd_sc_hd__clkbuf_1
X_4583_ _5140_/A VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__clkbuf_2
X_6322_ _7330_/A VGND VGND VPWR VPWR _7938_/A sky130_fd_sc_hd__buf_2
X_9041_ _9041_/A _9041_/B VGND VGND VPWR VPWR _9041_/Y sky130_fd_sc_hd__nor2_1
X_6253_ _7083_/A VGND VGND VPWR VPWR _7419_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5204_ _5204_/A VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__buf_2
X_6184_ _6182_/Y _6183_/X _6104_/C _6104_/Y VGND VGND VPWR VPWR _6207_/B sky130_fd_sc_hd__o211ai_2
XFILLER_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5135_ _5135_/A VGND VGND VPWR VPWR _5410_/A sky130_fd_sc_hd__clkbuf_2
X_5066_ _5164_/A _5064_/Y _5065_/X _4605_/A VGND VGND VPWR VPWR _5066_/X sky130_fd_sc_hd__a31o_1
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8825_ _8825_/A _8825_/B _8825_/C VGND VGND VPWR VPWR _8825_/Y sky130_fd_sc_hd__nand3_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8756_ _8756_/A _8756_/B VGND VGND VPWR VPWR _8757_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ _5968_/A _5968_/B _5968_/C VGND VGND VPWR VPWR _5976_/A sky130_fd_sc_hd__nand3_1
X_7707_ _7707_/A _7828_/A VGND VGND VPWR VPWR _7819_/C sky130_fd_sc_hd__nor2_1
X_4919_ _4943_/B VGND VGND VPWR VPWR _4920_/A sky130_fd_sc_hd__clkbuf_2
X_8687_ _8688_/B _8688_/C _8688_/A VGND VGND VPWR VPWR _8687_/Y sky130_fd_sc_hd__a21oi_1
X_5899_ _6014_/A _7367_/A _7367_/B _6169_/A VGND VGND VPWR VPWR _5903_/B sky130_fd_sc_hd__nand4_2
X_7638_ _8091_/D VGND VGND VPWR VPWR _8607_/D sky130_fd_sc_hd__buf_2
X_7569_ _7567_/X _7571_/A _7569_/C _7569_/D VGND VGND VPWR VPWR _7570_/B sky130_fd_sc_hd__and4b_1
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6940_ _6940_/A _6940_/B _6940_/C _6940_/D VGND VGND VPWR VPWR _6940_/Y sky130_fd_sc_hd__nor4_1
XFILLER_47_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6871_ _7419_/C VGND VGND VPWR VPWR _7923_/C sky130_fd_sc_hd__clkbuf_2
X_8610_ _8674_/A _8724_/A _8610_/C VGND VGND VPWR VPWR _8662_/B sky130_fd_sc_hd__and3_1
XFILLER_62_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _5818_/X _5940_/A _6031_/A _7506_/A VGND VGND VPWR VPWR _5870_/B sky130_fd_sc_hd__a22o_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8541_ _8664_/B _8542_/C _8239_/D _8664_/A VGND VGND VPWR VPWR _8543_/A sky130_fd_sc_hd__a22oi_1
X_5753_ _5484_/A _4875_/S _5752_/X _5749_/A VGND VGND VPWR VPWR _5754_/C sky130_fd_sc_hd__o22a_1
X_4704_ _4776_/A _4691_/A _4780_/A VGND VGND VPWR VPWR _4705_/B sky130_fd_sc_hd__a21oi_1
X_8472_ _8472_/A _8472_/B VGND VGND VPWR VPWR _8473_/B sky130_fd_sc_hd__nor2_1
X_5684_ _5450_/A _9097_/Q _4789_/A VGND VGND VPWR VPWR _5684_/Y sky130_fd_sc_hd__a21oi_1
X_7423_ _9213_/Q VGND VGND VPWR VPWR _7810_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4635_ _4635_/A VGND VGND VPWR VPWR _5402_/A sky130_fd_sc_hd__clkbuf_2
X_7354_ _7354_/A _7474_/A VGND VGND VPWR VPWR _7355_/B sky130_fd_sc_hd__and2_1
X_4566_ _4566_/A VGND VGND VPWR VPWR _4566_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6305_ _6302_/A _6302_/B _6304_/Y _6300_/B VGND VGND VPWR VPWR _6383_/A sky130_fd_sc_hd__a31oi_1
X_9024_ _8974_/Y _9002_/B _9009_/A VGND VGND VPWR VPWR _9027_/A sky130_fd_sc_hd__o21ai_1
X_7285_ _7285_/A _7285_/B VGND VGND VPWR VPWR _7287_/C sky130_fd_sc_hd__and2_1
X_6236_ _9173_/Q VGND VGND VPWR VPWR _7330_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6167_ _6097_/B _6100_/B _6097_/A VGND VGND VPWR VPWR _6268_/A sky130_fd_sc_hd__o21ba_1
XFILLER_84_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5118_ _9088_/Q VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__buf_2
X_6098_ _7129_/A VGND VGND VPWR VPWR _7988_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5049_ _4844_/X _5080_/B _5046_/B _5692_/S VGND VGND VPWR VPWR _5049_/X sky130_fd_sc_hd__a31o_1
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8808_ _8809_/A _8809_/B VGND VGND VPWR VPWR _8810_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8739_ _8816_/A _8798_/B VGND VGND VPWR VPWR _8741_/B sky130_fd_sc_hd__and2_1
XFILLER_68_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7070_ _7070_/A VGND VGND VPWR VPWR _7071_/C sky130_fd_sc_hd__inv_2
XFILLER_98_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6021_/A _6021_/B _6021_/C VGND VGND VPWR VPWR _6036_/C sky130_fd_sc_hd__and3_1
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7972_ _8102_/B _7972_/B VGND VGND VPWR VPWR _7974_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6923_ _6923_/A _6923_/B VGND VGND VPWR VPWR _6924_/B sky130_fd_sc_hd__nor2_1
X_6854_ _7824_/B VGND VGND VPWR VPWR _8052_/B sky130_fd_sc_hd__buf_2
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6785_ _9196_/Q VGND VGND VPWR VPWR _7259_/A sky130_fd_sc_hd__buf_2
X_5805_ _9196_/Q VGND VGND VPWR VPWR _7367_/A sky130_fd_sc_hd__buf_2
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8524_ _8525_/A _8525_/B _8525_/C VGND VGND VPWR VPWR _8624_/A sky130_fd_sc_hd__a21oi_1
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5736_ _4641_/A _5735_/X _5736_/S VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__mux2_1
X_8455_ _8639_/A _8975_/A VGND VGND VPWR VPWR _8456_/B sky130_fd_sc_hd__nand2_1
X_5667_ _5432_/A _5712_/S _5666_/X VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7406_ _7406_/A _7552_/A _7552_/B VGND VGND VPWR VPWR _7408_/B sky130_fd_sc_hd__and3_1
X_4618_ _9108_/Q VGND VGND VPWR VPWR _5739_/S sky130_fd_sc_hd__inv_2
X_8386_ _8466_/A _8542_/A _8464_/B _8664_/B VGND VGND VPWR VPWR _8387_/B sky130_fd_sc_hd__and4_1
X_5598_ _5433_/A _4799_/A _5596_/X _5597_/Y VGND VGND VPWR VPWR _5598_/X sky130_fd_sc_hd__a22o_1
X_7337_ _7338_/A _7338_/B VGND VGND VPWR VPWR _7339_/A sky130_fd_sc_hd__nor2_1
X_4549_ _5129_/A VGND VGND VPWR VPWR _4550_/A sky130_fd_sc_hd__buf_2
X_7268_ _7377_/B _7377_/C _7377_/A VGND VGND VPWR VPWR _7268_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9007_ _8982_/A _8982_/B _9006_/Y VGND VGND VPWR VPWR _9008_/B sky130_fd_sc_hd__a21boi_1
X_6219_ _6302_/B _6219_/B VGND VGND VPWR VPWR _6220_/A sky130_fd_sc_hd__and2_1
X_7199_ _7199_/A _7307_/A _7822_/C _7307_/D VGND VGND VPWR VPWR _7200_/B sky130_fd_sc_hd__and4_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6570_ _6968_/A _7962_/B VGND VGND VPWR VPWR _6571_/B sky130_fd_sc_hd__nand2_1
X_5521_ _5213_/X _5420_/X _5519_/X _5520_/Y _5227_/X VGND VGND VPWR VPWR _5521_/X
+ sky130_fd_sc_hd__a221o_1
X_8240_ _8240_/A _8240_/B VGND VGND VPWR VPWR _8242_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5452_ _5315_/X _5187_/X _5448_/X _5451_/Y VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__a22o_1
X_8171_ _8082_/B _8107_/A _8266_/A _8169_/Y VGND VGND VPWR VPWR _8171_/X sky130_fd_sc_hd__a211o_1
X_5383_ _5382_/X _5273_/X _5170_/X VGND VGND VPWR VPWR _5383_/Y sky130_fd_sc_hd__a21oi_1
X_7122_ _7122_/A _7122_/B VGND VGND VPWR VPWR _7124_/A sky130_fd_sc_hd__xnor2_1
X_7053_ _7053_/A _7053_/B _7053_/C VGND VGND VPWR VPWR _7053_/Y sky130_fd_sc_hd__nor3_2
XFILLER_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6004_ _6447_/A _9167_/Q _6232_/A _6055_/A VGND VGND VPWR VPWR _6007_/C sky130_fd_sc_hd__a22o_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _7832_/B _7837_/C _7952_/X _8029_/A VGND VGND VPWR VPWR _8029_/B sky130_fd_sc_hd__a211oi_2
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7886_ _7984_/A _7997_/A _7885_/X VGND VGND VPWR VPWR _7888_/A sky130_fd_sc_hd__o21ai_1
X_6906_ _7986_/A _7938_/A _7938_/B _7869_/A VGND VGND VPWR VPWR _6908_/A sky130_fd_sc_hd__a22oi_1
XFILLER_23_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6837_ _6837_/A _6837_/B VGND VGND VPWR VPWR _6945_/A sky130_fd_sc_hd__xor2_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8507_ _8513_/A _8513_/B VGND VGND VPWR VPWR _8580_/A sky130_fd_sc_hd__xnor2_2
X_6768_ _6767_/A _6767_/B _6767_/C VGND VGND VPWR VPWR _6879_/A sky130_fd_sc_hd__a21oi_4
X_5719_ _5714_/S _5765_/B _4891_/X _5718_/X VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__a211o_1
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6699_ _9207_/Q VGND VGND VPWR VPWR _7849_/B sky130_fd_sc_hd__buf_2
X_8438_ _8438_/A _8438_/B _8841_/A _8842_/B VGND VGND VPWR VPWR _8439_/B sky130_fd_sc_hd__and4_1
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8369_ _8452_/A _8379_/A _8842_/A _8733_/D VGND VGND VPWR VPWR _8370_/B sky130_fd_sc_hd__and4_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 A[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7740_ _7740_/A _7740_/B _7740_/C VGND VGND VPWR VPWR _7745_/B sky130_fd_sc_hd__nand3_1
XFILLER_91_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4952_ _5158_/A _4949_/Y _4951_/X VGND VGND VPWR VPWR _4952_/X sky130_fd_sc_hd__o21a_1
X_4883_ _5403_/A VGND VGND VPWR VPWR _4883_/X sky130_fd_sc_hd__clkbuf_2
X_7671_ _7672_/A _7672_/B VGND VGND VPWR VPWR _7795_/A sky130_fd_sc_hd__or2_1
X_6622_ _6622_/A _6622_/B VGND VGND VPWR VPWR _6637_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6553_ _6553_/A _6553_/B VGND VGND VPWR VPWR _6655_/A sky130_fd_sc_hd__xnor2_2
X_6484_ _6646_/A _6484_/B VGND VGND VPWR VPWR _6553_/A sky130_fd_sc_hd__and2_1
X_5504_ _5628_/A VGND VGND VPWR VPWR _5603_/S sky130_fd_sc_hd__clkbuf_2
X_8223_ _8223_/A _8223_/B _8223_/C VGND VGND VPWR VPWR _8224_/B sky130_fd_sc_hd__nor3_1
X_5435_ _5558_/A _5248_/A _4580_/X _5507_/A _5434_/Y VGND VGND VPWR VPWR _5435_/X
+ sky130_fd_sc_hd__o221a_1
X_8154_ _8154_/A _8154_/B VGND VGND VPWR VPWR _8154_/X sky130_fd_sc_hd__and2_1
X_5366_ _5511_/A VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__clkbuf_2
X_8085_ _8516_/A _8466_/A _8150_/C _8086_/A VGND VGND VPWR VPWR _8087_/A sky130_fd_sc_hd__a22oi_1
X_5297_ _5382_/A _5179_/X _4641_/A VGND VGND VPWR VPWR _5297_/Y sky130_fd_sc_hd__a21oi_1
X_7105_ _7104_/A _7104_/B _7104_/C VGND VGND VPWR VPWR _7281_/B sky130_fd_sc_hd__a21oi_2
X_7036_ _7694_/B _6493_/C _7728_/D _7146_/A VGND VGND VPWR VPWR _7038_/A sky130_fd_sc_hd__a22oi_1
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8987_ _8932_/A _8932_/B _8936_/B VGND VGND VPWR VPWR _8988_/B sky130_fd_sc_hd__a21oi_2
XFILLER_82_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _7938_/A _7938_/B _7938_/C _8050_/D VGND VGND VPWR VPWR _8056_/A sky130_fd_sc_hd__and4_1
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7869_ _7869_/A _8154_/B VGND VGND VPWR VPWR _8068_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5220_ _4585_/A _5316_/A _5218_/Y _5219_/X VGND VGND VPWR VPWR _5220_/X sky130_fd_sc_hd__a211o_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5151_ _5151_/A VGND VGND VPWR VPWR _5151_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5082_ _5048_/Y _5049_/X _5078_/X _5081_/X VGND VGND VPWR VPWR _5082_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8910_ _8959_/A _8959_/B VGND VGND VPWR VPWR _8957_/B sky130_fd_sc_hd__xnor2_2
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8841_ _8841_/A VGND VGND VPWR VPWR _8989_/A sky130_fd_sc_hd__buf_2
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8772_ _8772_/A _8772_/B VGND VGND VPWR VPWR _8772_/X sky130_fd_sc_hd__and2_1
X_5984_ _7349_/A VGND VGND VPWR VPWR _6172_/A sky130_fd_sc_hd__clkbuf_2
X_7723_ _7724_/B _7724_/C _7724_/A VGND VGND VPWR VPWR _7725_/A sky130_fd_sc_hd__a21oi_1
X_4935_ _4935_/A VGND VGND VPWR VPWR _5146_/A sky130_fd_sc_hd__buf_2
XANTENNA_11 _9154_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7654_ _7764_/A _7764_/B VGND VGND VPWR VPWR _7776_/B sky130_fd_sc_hd__xor2_2
XANTENNA_22 _9137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4866_ _4866_/A _4960_/B VGND VGND VPWR VPWR _4915_/A sky130_fd_sc_hd__nor2_2
X_7585_ _7925_/A _8185_/A _7586_/C VGND VGND VPWR VPWR _7587_/A sky130_fd_sc_hd__a21oi_1
X_6605_ _6760_/A _6680_/B _7327_/A _6680_/A VGND VGND VPWR VPWR _6606_/B sky130_fd_sc_hd__a22oi_2
XANTENNA_33 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _9071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _9195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4769_/B _4796_/X _5691_/S VGND VGND VPWR VPWR _4797_/X sky130_fd_sc_hd__mux2_1
X_6536_ _6536_/A _6536_/B VGND VGND VPWR VPWR _6537_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6467_ _6551_/B _6465_/X _6372_/C _6466_/Y VGND VGND VPWR VPWR _6469_/A sky130_fd_sc_hd__a211oi_1
X_9186_ _9222_/CLK _9186_/D VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
X_8206_ _8060_/B _8063_/B _8203_/X _8318_/A VGND VGND VPWR VPWR _8318_/B sky130_fd_sc_hd__a211oi_2
X_5418_ _5177_/X _5120_/A _5416_/X _5417_/Y _4545_/A VGND VGND VPWR VPWR _5418_/X
+ sky130_fd_sc_hd__a221o_1
X_6398_ _7189_/C _6828_/A _7847_/A _7459_/D VGND VGND VPWR VPWR _6483_/A sky130_fd_sc_hd__and4_2
X_8137_ _8137_/A _8587_/B VGND VGND VPWR VPWR _8138_/B sky130_fd_sc_hd__nand2_1
X_5349_ _5213_/X _5184_/X _5347_/X _5348_/Y _5227_/X VGND VGND VPWR VPWR _5349_/X
+ sky130_fd_sc_hd__a221o_1
X_8068_ _8068_/A _8257_/C VGND VGND VPWR VPWR _8078_/A sky130_fd_sc_hd__nor2_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7019_ _7131_/A _7019_/B _7019_/C _9175_/Q VGND VGND VPWR VPWR _7020_/B sky130_fd_sc_hd__and4_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4875_/S _4717_/X _4719_/X VGND VGND VPWR VPWR _4720_/X sky130_fd_sc_hd__a21o_1
X_4651_ _9108_/Q VGND VGND VPWR VPWR _5103_/A sky130_fd_sc_hd__clkbuf_2
Xinput31 A[8] VGND VGND VPWR VPWR _9170_/D sky130_fd_sc_hd__clkbuf_1
Xinput20 A[27] VGND VGND VPWR VPWR _9189_/D sky130_fd_sc_hd__clkbuf_1
X_7370_ _7261_/A _7260_/A _7260_/B VGND VGND VPWR VPWR _7371_/B sky130_fd_sc_hd__o21ba_1
Xinput53 B[28] VGND VGND VPWR VPWR _9221_/D sky130_fd_sc_hd__clkbuf_2
Xinput42 B[18] VGND VGND VPWR VPWR _9211_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 B[9] VGND VGND VPWR VPWR _9202_/D sky130_fd_sc_hd__clkbuf_1
X_4582_ _4582_/A VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__clkbuf_2
X_6321_ _6321_/A _6321_/B VGND VGND VPWR VPWR _6434_/A sky130_fd_sc_hd__xnor2_4
X_9040_ _9040_/A _9040_/B VGND VGND VPWR VPWR _9110_/D sky130_fd_sc_hd__xnor2_1
X_6252_ _7187_/A _6607_/B VGND VGND VPWR VPWR _6259_/A sky130_fd_sc_hd__nand2_1
X_5203_ _5511_/A VGND VGND VPWR VPWR _5204_/A sky130_fd_sc_hd__clkbuf_2
X_6183_ _6264_/A _6264_/B _6264_/C VGND VGND VPWR VPWR _6183_/X sky130_fd_sc_hd__and3_1
X_5134_ _5248_/A VGND VGND VPWR VPWR _5532_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5065_ _5065_/A _5067_/B _5072_/A VGND VGND VPWR VPWR _5065_/X sky130_fd_sc_hd__or3_1
XFILLER_65_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8824_ _8825_/A _8825_/B _8825_/C VGND VGND VPWR VPWR _8826_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8755_ _8755_/A _8755_/B VGND VGND VPWR VPWR _8757_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5967_ _5903_/A _5903_/C _5903_/B VGND VGND VPWR VPWR _5968_/C sky130_fd_sc_hd__a21bo_1
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8686_ _8686_/A _8686_/B _8745_/A VGND VGND VPWR VPWR _8688_/C sky130_fd_sc_hd__or3_1
X_7706_ _7706_/A _7706_/B _7706_/C _7706_/D VGND VGND VPWR VPWR _7828_/A sky130_fd_sc_hd__and4_1
X_4918_ _5740_/S VGND VGND VPWR VPWR _5696_/S sky130_fd_sc_hd__buf_2
X_7637_ _7637_/A _7726_/A VGND VGND VPWR VPWR _7657_/A sky130_fd_sc_hd__xnor2_2
X_5898_ _5862_/X _5898_/B _5898_/C VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__and3b_1
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4849_ _4849_/A VGND VGND VPWR VPWR _5144_/A sky130_fd_sc_hd__clkbuf_2
X_7568_ _7569_/C _7810_/B _7566_/Y _7567_/X VGND VGND VPWR VPWR _7570_/A sky130_fd_sc_hd__o2bb2a_1
X_7499_ _7499_/A VGND VGND VPWR VPWR _7880_/A sky130_fd_sc_hd__clkbuf_2
X_6519_ _7810_/C _7485_/A _6521_/C VGND VGND VPWR VPWR _6565_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9169_ _9224_/CLK _9169_/D VGND VGND VPWR VPWR _9169_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6870_ _9211_/Q VGND VGND VPWR VPWR _7419_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5821_ _6139_/A VGND VGND VPWR VPWR _7506_/A sky130_fd_sc_hd__buf_2
X_8540_ _8439_/A _8442_/B _8439_/B VGND VGND VPWR VPWR _8547_/A sky130_fd_sc_hd__o21ba_1
X_5752_ _5364_/A _5621_/X _4636_/A _4637_/A _5751_/Y VGND VGND VPWR VPWR _5752_/X
+ sky130_fd_sc_hd__o32a_1
X_4703_ _5732_/S VGND VGND VPWR VPWR _4875_/S sky130_fd_sc_hd__clkbuf_2
X_8471_ _8470_/A _8470_/B _8470_/C VGND VGND VPWR VPWR _8472_/B sky130_fd_sc_hd__o21a_1
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5683_ _9091_/Q _4861_/A _5682_/X _9097_/Q VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__a211o_1
X_7422_ _7422_/A _7422_/B VGND VGND VPWR VPWR _7425_/A sky130_fd_sc_hd__nor2_1
X_4634_ _4634_/A VGND VGND VPWR VPWR _4635_/A sky130_fd_sc_hd__clkbuf_2
X_7353_ _7352_/A _7352_/B _7352_/C VGND VGND VPWR VPWR _7474_/A sky130_fd_sc_hd__o21ai_2
X_4565_ _4786_/S VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6304_ _6304_/A _6304_/B _6304_/C VGND VGND VPWR VPWR _6304_/Y sky130_fd_sc_hd__nand3_1
X_9023_ _9023_/A _9017_/A VGND VGND VPWR VPWR _9035_/B sky130_fd_sc_hd__or2b_1
X_7284_ _7284_/A _7284_/B _7284_/C VGND VGND VPWR VPWR _7285_/B sky130_fd_sc_hd__nand3_1
XFILLER_103_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6235_ _6235_/A VGND VGND VPWR VPWR _6998_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A _6166_/B _6166_/C VGND VGND VPWR VPWR _6264_/C sky130_fd_sc_hd__nand3_2
XFILLER_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5117_ _5117_/A VGND VGND VPWR VPWR _5117_/X sky130_fd_sc_hd__buf_2
X_6097_ _6097_/A _6097_/B VGND VGND VPWR VPWR _6100_/A sky130_fd_sc_hd__nor2_1
X_5048_ _4844_/X _5046_/B _5040_/A VGND VGND VPWR VPWR _5048_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8807_ _8863_/A _8807_/B VGND VGND VPWR VPWR _8809_/B sky130_fd_sc_hd__xor2_1
XFILLER_53_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6999_ _7259_/D VGND VGND VPWR VPWR _7988_/B sky130_fd_sc_hd__buf_2
X_8738_ _8738_/A _8811_/A VGND VGND VPWR VPWR _8741_/A sky130_fd_sc_hd__xnor2_1
XFILLER_80_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A VGND VGND VPWR VPWR _9214_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8669_ _8668_/A _8668_/B _8668_/C VGND VGND VPWR VPWR _8670_/B sky130_fd_sc_hd__o21a_1
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6020_ _6021_/A _6021_/B _6021_/C VGND VGND VPWR VPWR _6036_/B sky130_fd_sc_hd__a21oi_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7971_ _7853_/A _7855_/B _7853_/B VGND VGND VPWR VPWR _7972_/B sky130_fd_sc_hd__o21ba_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6922_ _7419_/B _6922_/B _7728_/B _7728_/D VGND VGND VPWR VPWR _6923_/B sky130_fd_sc_hd__and4_1
XFILLER_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6853_ _6853_/A VGND VGND VPWR VPWR _6882_/A sky130_fd_sc_hd__inv_2
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5804_ _9163_/Q VGND VGND VPWR VPWR _5940_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6784_ _7257_/A _7852_/C VGND VGND VPWR VPWR _6791_/A sky130_fd_sc_hd__nand2_1
X_8523_ _8523_/A _8523_/B VGND VGND VPWR VPWR _8525_/C sky130_fd_sc_hd__xnor2_1
X_5735_ _4923_/A _5734_/X _5735_/S VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__mux2_1
X_8454_ _8794_/B VGND VGND VPWR VPWR _8975_/A sky130_fd_sc_hd__clkbuf_2
X_5666_ _4634_/A _5071_/A _5664_/X _5665_/Y _4721_/A VGND VGND VPWR VPWR _5666_/X
+ sky130_fd_sc_hd__a221o_1
X_4617_ _5632_/A _4613_/X _5676_/A VGND VGND VPWR VPWR _4617_/X sky130_fd_sc_hd__o21a_1
X_7405_ _7405_/A _7547_/B VGND VGND VPWR VPWR _7408_/A sky130_fd_sc_hd__xnor2_2
X_8385_ _8664_/A _8675_/A _8831_/A _8595_/A VGND VGND VPWR VPWR _8387_/A sky130_fd_sc_hd__a22oi_1
X_5597_ _4566_/X _5271_/A _5181_/A VGND VGND VPWR VPWR _5597_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7336_ _7476_/B _7336_/B VGND VGND VPWR VPWR _7338_/B sky130_fd_sc_hd__xnor2_1
X_4548_ _4548_/A VGND VGND VPWR VPWR _5129_/A sky130_fd_sc_hd__clkbuf_2
X_7267_ _7377_/A _7377_/B _7377_/C VGND VGND VPWR VPWR _7267_/X sky130_fd_sc_hd__and3_1
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9006_ _9006_/A _9006_/B VGND VGND VPWR VPWR _9006_/Y sky130_fd_sc_hd__xnor2_1
X_6218_ _6218_/A _6218_/B _6218_/C VGND VGND VPWR VPWR _6219_/B sky130_fd_sc_hd__nand3_1
X_7198_ _6572_/B _6825_/C _7706_/D _6500_/B VGND VGND VPWR VPWR _7200_/A sky130_fd_sc_hd__a22oi_1
X_6149_ _9172_/Q VGND VGND VPWR VPWR _7327_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5520_ _4717_/S _5119_/A _5213_/A VGND VGND VPWR VPWR _5520_/Y sky130_fd_sc_hd__a21oi_1
X_5451_ _5450_/X _5276_/X _5105_/A VGND VGND VPWR VPWR _5451_/Y sky130_fd_sc_hd__a21oi_1
X_8170_ _8266_/A _8169_/Y _8082_/B _8107_/A VGND VGND VPWR VPWR _8172_/A sky130_fd_sc_hd__o211a_1
X_5382_ _5382_/A VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__clkbuf_2
X_7121_ _7121_/A _7121_/B VGND VGND VPWR VPWR _7122_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7052_ _7053_/B _7053_/C _7053_/A VGND VGND VPWR VPWR _7052_/X sky130_fd_sc_hd__o21a_1
X_6003_ _6139_/A _7259_/B _6256_/A _6232_/A VGND VGND VPWR VPWR _6007_/B sky130_fd_sc_hd__nand4_2
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7954_ _7952_/X _8029_/A _7832_/B _7837_/C VGND VGND VPWR VPWR _7956_/A sky130_fd_sc_hd__o211a_1
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _7988_/A _7602_/A VGND VGND VPWR VPWR _6909_/A sky130_fd_sc_hd__nand2_1
X_7885_ _7880_/A _8831_/B _8780_/B _7766_/A VGND VGND VPWR VPWR _7885_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _6836_/A _6835_/X VGND VGND VPWR VPWR _6837_/B sky130_fd_sc_hd__or2b_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6767_ _6767_/A _6767_/B _6767_/C VGND VGND VPWR VPWR _6772_/B sky130_fd_sc_hd__and3_1
X_8506_ _8415_/A _9025_/B _8416_/A _8414_/B VGND VGND VPWR VPWR _8513_/B sky130_fd_sc_hd__a31oi_4
X_5718_ _5713_/S _5765_/C _5716_/Y _5717_/X _5281_/S VGND VGND VPWR VPWR _5718_/X
+ sky130_fd_sc_hd__o221a_1
X_6698_ _6696_/X _6698_/B VGND VGND VPWR VPWR _6701_/A sky130_fd_sc_hd__and2b_1
X_8437_ _8438_/B _8844_/B _8842_/B _8438_/A VGND VGND VPWR VPWR _8439_/A sky130_fd_sc_hd__a22oi_1
X_5649_ _5509_/A _4999_/X _5765_/C _5648_/X VGND VGND VPWR VPWR _5649_/Y sky130_fd_sc_hd__o211ai_1
X_8368_ _8595_/C VGND VGND VPWR VPWR _8842_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7319_ _7319_/A _7319_/B _7319_/C VGND VGND VPWR VPWR _7319_/X sky130_fd_sc_hd__and3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8299_ _8299_/A _8299_/B _8299_/C VGND VGND VPWR VPWR _8300_/B sky130_fd_sc_hd__nor3_1
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 A[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4951_ _5729_/S _4951_/B _5052_/A VGND VGND VPWR VPWR _4951_/X sky130_fd_sc_hd__or3_1
X_4882_ _5606_/A _4882_/B VGND VGND VPWR VPWR _4882_/Y sky130_fd_sc_hd__nand2_1
X_7670_ _7670_/A _7793_/A VGND VGND VPWR VPWR _7672_/B sky130_fd_sc_hd__and2_1
X_6621_ _6548_/C _6550_/A _6618_/X _6619_/Y VGND VGND VPWR VPWR _6640_/C sky130_fd_sc_hd__o211ai_1
X_6552_ _6643_/A _6643_/B VGND VGND VPWR VPWR _6553_/B sky130_fd_sc_hd__xnor2_1
X_6483_ _6483_/A _6483_/B _6483_/C VGND VGND VPWR VPWR _6484_/B sky130_fd_sc_hd__or3_1
X_5503_ _5433_/X _5502_/X _5553_/S VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
X_8222_ _8223_/B _8223_/C _8223_/A VGND VGND VPWR VPWR _8224_/A sky130_fd_sc_hd__o21a_1
X_5434_ _5404_/A _5146_/X _4847_/X VGND VGND VPWR VPWR _5434_/Y sky130_fd_sc_hd__a21oi_1
X_8153_ _8153_/A _8153_/B VGND VGND VPWR VPWR _8162_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5365_ _5365_/A VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__clkbuf_2
X_7104_ _7104_/A _7104_/B _7104_/C VGND VGND VPWR VPWR _7104_/X sky130_fd_sc_hd__and3_1
XFILLER_101_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8084_ _8084_/A VGND VGND VPWR VPWR _8516_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5296_ _5367_/A _5581_/A _5294_/X _5295_/Y _5132_/A VGND VGND VPWR VPWR _5296_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7035_ _7309_/A _9207_/Q VGND VGND VPWR VPWR _7039_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8986_ _9006_/B _8986_/B VGND VGND VPWR VPWR _8992_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7937_ _7604_/B _8050_/C _8720_/A _7730_/A VGND VGND VPWR VPWR _7939_/A sky130_fd_sc_hd__a22oi_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _7747_/X _8733_/A _7759_/A _7754_/Y VGND VGND VPWR VPWR _7878_/A sky130_fd_sc_hd__a31o_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ _7562_/A _7849_/B _6698_/B _6696_/X VGND VGND VPWR VPWR _6830_/A sky130_fd_sc_hd__a31o_2
XFILLER_23_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7799_ _7799_/A _7799_/B VGND VGND VPWR VPWR _7903_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5150_ _9071_/Q VGND VGND VPWR VPWR _5150_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5081_ _4878_/A _5079_/Y _5080_/X _5125_/A VGND VGND VPWR VPWR _5081_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_8840_ _8840_/A _8904_/A VGND VGND VPWR VPWR _8855_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8771_ _8771_/A _8771_/B VGND VGND VPWR VPWR _8772_/B sky130_fd_sc_hd__nor2_1
X_5983_ _6825_/B _6257_/C _6424_/D _6031_/A VGND VGND VPWR VPWR _5986_/A sky130_fd_sc_hd__a22oi_2
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7722_ _7592_/A _7592_/B _7594_/Y VGND VGND VPWR VPWR _7724_/A sky130_fd_sc_hd__o21bai_1
X_4934_ _5656_/B _4932_/X _4933_/Y _4783_/X VGND VGND VPWR VPWR _4934_/X sky130_fd_sc_hd__a31o_1
X_7653_ _7653_/A _7772_/A VGND VGND VPWR VPWR _7764_/B sky130_fd_sc_hd__nor2_1
XANTENNA_12 _9155_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _5424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ _5054_/S _4950_/A VGND VGND VPWR VPWR _5080_/A sky130_fd_sc_hd__nor2_1
X_7584_ _7584_/A _7712_/A VGND VGND VPWR VPWR _7586_/C sky130_fd_sc_hd__nor2_1
X_6604_ _7131_/A _9170_/Q _7347_/A _9171_/Q VGND VGND VPWR VPWR _6606_/A sky130_fd_sc_hd__and4_1
XANTENNA_34 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 _9198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _9140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4796_ _4773_/Y _4795_/Y _5734_/S VGND VGND VPWR VPWR _4796_/X sky130_fd_sc_hd__mux2_1
X_6535_ _6223_/A _7455_/A _7129_/B _6223_/B VGND VGND VPWR VPWR _6536_/B sky130_fd_sc_hd__a22oi_2
X_8205_ _8203_/X _8318_/A _8060_/B _8063_/B VGND VGND VPWR VPWR _8207_/A sky130_fd_sc_hd__o211a_1
X_6466_ _6466_/A VGND VGND VPWR VPWR _6466_/Y sky130_fd_sc_hd__inv_2
X_6397_ _7728_/D VGND VGND VPWR VPWR _7459_/D sky130_fd_sc_hd__buf_2
X_5417_ _5385_/X _5194_/X _4656_/A VGND VGND VPWR VPWR _5417_/Y sky130_fd_sc_hd__a21oi_1
X_9185_ _9199_/CLK _9185_/D VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
X_8136_ _7747_/X _8831_/B _8780_/B _8069_/A VGND VGND VPWR VPWR _8139_/A sky130_fd_sc_hd__a22o_1
X_5348_ _4717_/S _5630_/A _4605_/A VGND VGND VPWR VPWR _5348_/Y sky130_fd_sc_hd__a21oi_1
X_8067_ _7948_/B _7951_/B _8064_/X _8217_/A VGND VGND VPWR VPWR _8217_/B sky130_fd_sc_hd__a211oi_2
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7018_ _5985_/D _7019_/C _7131_/C _6172_/A VGND VGND VPWR VPWR _7020_/A sky130_fd_sc_hd__a22oi_1
XFILLER_75_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5279_ _5276_/X _5278_/X _5105_/A VGND VGND VPWR VPWR _5279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8969_ _8920_/A _8920_/B _8967_/Y _8881_/X _8968_/X VGND VGND VPWR VPWR _8970_/A
+ sky130_fd_sc_hd__a221oi_1
XFILLER_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _4650_/A VGND VGND VPWR VPWR _5339_/A sky130_fd_sc_hd__buf_2
Xinput21 A[28] VGND VGND VPWR VPWR _9190_/D sky130_fd_sc_hd__clkbuf_1
Xinput10 A[18] VGND VGND VPWR VPWR _9180_/D sky130_fd_sc_hd__clkbuf_1
Xinput32 A[9] VGND VGND VPWR VPWR _9171_/D sky130_fd_sc_hd__clkbuf_1
Xinput54 B[29] VGND VGND VPWR VPWR _9222_/D sky130_fd_sc_hd__clkbuf_1
Xinput43 B[19] VGND VGND VPWR VPWR _9212_/D sky130_fd_sc_hd__clkbuf_1
X_6320_ _6320_/A _6320_/B VGND VGND VPWR VPWR _6321_/B sky130_fd_sc_hd__nor2_2
X_4581_ _9095_/Q VGND VGND VPWR VPWR _4582_/A sky130_fd_sc_hd__clkbuf_2
X_6251_ _6251_/A VGND VGND VPWR VPWR _7187_/A sky130_fd_sc_hd__clkbuf_2
X_5202_ _5365_/A VGND VGND VPWR VPWR _5202_/X sky130_fd_sc_hd__buf_2
X_6182_ _6264_/B _6264_/C _6264_/A VGND VGND VPWR VPWR _6182_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5133_ _9078_/Q VGND VGND VPWR VPWR _5248_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5064_ _5065_/A _5072_/A _5074_/B VGND VGND VPWR VPWR _5064_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8823_ _8829_/A _8829_/B VGND VGND VPWR VPWR _8825_/C sky130_fd_sc_hd__xnor2_1
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8754_ _8753_/A _8753_/B _8752_/Y VGND VGND VPWR VPWR _8755_/B sky130_fd_sc_hd__o21ba_1
XFILLER_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5966_ _5965_/A _5965_/C _5965_/B VGND VGND VPWR VPWR _5968_/B sky130_fd_sc_hd__o21ai_1
X_8685_ _8686_/B _8745_/A _8686_/A VGND VGND VPWR VPWR _8688_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7705_ _7457_/A _7938_/C _8050_/D _7583_/B VGND VGND VPWR VPWR _7707_/A sky130_fd_sc_hd__a22oi_1
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5897_ _5897_/A VGND VGND VPWR VPWR _5951_/A sky130_fd_sc_hd__inv_2
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4917_ _9109_/Q VGND VGND VPWR VPWR _5740_/S sky130_fd_sc_hd__clkinv_2
X_7636_ _7636_/A _7740_/A VGND VGND VPWR VPWR _7726_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4848_ _4940_/A VGND VGND VPWR VPWR _4849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7567_ _7696_/C _7694_/A _7923_/C _7923_/D VGND VGND VPWR VPWR _7567_/X sky130_fd_sc_hd__and4_1
X_4779_ _9093_/Q _9092_/Q VGND VGND VPWR VPWR _4935_/A sky130_fd_sc_hd__nor2_1
X_7498_ _7766_/A _8156_/C VGND VGND VPWR VPWR _7643_/A sky130_fd_sc_hd__nand2_1
X_6518_ _6611_/A _6518_/B VGND VGND VPWR VPWR _6521_/C sky130_fd_sc_hd__nor2_1
X_6449_ _7152_/D VGND VGND VPWR VPWR _7822_/B sky130_fd_sc_hd__buf_2
XFILLER_79_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9168_ _9220_/CLK _9168_/D VGND VGND VPWR VPWR _9168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8119_ _8012_/A _8012_/B _8118_/X VGND VGND VPWR VPWR _8120_/B sky130_fd_sc_hd__a21bo_1
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9099_ _9221_/CLK _9099_/D VGND VGND VPWR VPWR _9099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5820_ _9196_/Q VGND VGND VPWR VPWR _6139_/A sky130_fd_sc_hd__clkbuf_2
X_5751_ _4573_/X _5621_/X _4635_/A _4560_/A VGND VGND VPWR VPWR _5751_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8470_ _8470_/A _8470_/B _8470_/C VGND VGND VPWR VPWR _8472_/A sky130_fd_sc_hd__nor3_1
X_4702_ _9101_/Q VGND VGND VPWR VPWR _5732_/S sky130_fd_sc_hd__inv_2
X_7421_ _7419_/X _7696_/B _7421_/C _7421_/D VGND VGND VPWR VPWR _7422_/B sky130_fd_sc_hd__and4b_1
X_5682_ _9090_/Q _4857_/A _5680_/X _5681_/X _5727_/S VGND VGND VPWR VPWR _5682_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ _5368_/A VGND VGND VPWR VPWR _4634_/A sky130_fd_sc_hd__clkbuf_2
X_7352_ _7352_/A _7352_/B _7352_/C VGND VGND VPWR VPWR _7354_/A sky130_fd_sc_hd__or3_1
X_4564_ _5727_/S VGND VGND VPWR VPWR _4786_/S sky130_fd_sc_hd__buf_2
X_6303_ _6303_/A _6303_/B VGND VGND VPWR VPWR _9078_/D sky130_fd_sc_hd__xnor2_1
X_7283_ _7284_/B _7284_/C _7284_/A VGND VGND VPWR VPWR _7285_/A sky130_fd_sc_hd__a21o_1
X_9022_ _9022_/A _9022_/B VGND VGND VPWR VPWR _9109_/D sky130_fd_sc_hd__xor2_1
X_6234_ _7146_/A _6775_/A VGND VGND VPWR VPWR _6335_/A sky130_fd_sc_hd__nand2_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6166_/A _6166_/B _6166_/C VGND VGND VPWR VPWR _6264_/B sky130_fd_sc_hd__a21o_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _7081_/A _7869_/A _7986_/A _6361_/B VGND VGND VPWR VPWR _6097_/B sky130_fd_sc_hd__a22oi_2
X_5116_ _5116_/A VGND VGND VPWR VPWR _5117_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5047_ _5040_/A _5046_/B _5181_/A VGND VGND VPWR VPWR _5047_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6998_ _6998_/A _6998_/B _7347_/B _7259_/D VGND VGND VPWR VPWR _7134_/A sky130_fd_sc_hd__and4_1
X_8806_ _8806_/A _8806_/B VGND VGND VPWR VPWR _8807_/B sky130_fd_sc_hd__nand2_1
X_8737_ _8678_/A _8680_/B _8678_/B VGND VGND VPWR VPWR _8811_/A sky130_fd_sc_hd__o21ba_1
XFILLER_80_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5949_ _9059_/A _9062_/A VGND VGND VPWR VPWR _9060_/B sky130_fd_sc_hd__and2_1
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8668_ _8668_/A _8668_/B _8668_/C VGND VGND VPWR VPWR _8670_/A sky130_fd_sc_hd__nor3_1
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7619_ _7473_/A _7473_/B _7618_/X VGND VGND VPWR VPWR _7621_/A sky130_fd_sc_hd__a21o_1
X_8599_ _8527_/A _8794_/B _8532_/D _8530_/X VGND VGND VPWR VPWR _8600_/B sky130_fd_sc_hd__a31o_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7970_ _7970_/A _7970_/B VGND VGND VPWR VPWR _8102_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6921_ _7694_/A _7604_/C _7847_/C _7309_/A VGND VGND VPWR VPWR _6923_/A sky130_fd_sc_hd__a22oi_1
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6852_ _6837_/A _6836_/A _6835_/X VGND VGND VPWR VPWR _6949_/A sky130_fd_sc_hd__o21a_2
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5803_ _7293_/A _7257_/A VGND VGND VPWR VPWR _5812_/A sky130_fd_sc_hd__nand2_2
X_8522_ _8522_/A _8522_/B VGND VGND VPWR VPWR _8523_/B sky130_fd_sc_hd__nor2_1
X_6783_ _7348_/B VGND VGND VPWR VPWR _7852_/C sky130_fd_sc_hd__clkbuf_2
X_5734_ _4716_/A _5733_/X _5734_/S VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__mux2_1
X_8453_ _8597_/B VGND VGND VPWR VPWR _8794_/B sky130_fd_sc_hd__clkbuf_2
X_5665_ _5618_/X _5213_/A _5227_/A VGND VGND VPWR VPWR _5665_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8384_ _8542_/B VGND VGND VPWR VPWR _8831_/A sky130_fd_sc_hd__clkbuf_2
X_4616_ _5354_/S VGND VGND VPWR VPWR _5676_/A sky130_fd_sc_hd__clkbuf_2
X_7404_ _7404_/A _7411_/A VGND VGND VPWR VPWR _7547_/B sky130_fd_sc_hd__nor2_1
X_7335_ _7335_/A _7342_/A VGND VGND VPWR VPWR _7336_/B sky130_fd_sc_hd__nor2_1
X_5596_ _4587_/X _5175_/A _5594_/X _5595_/Y _5125_/A VGND VGND VPWR VPWR _5596_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _4721_/A VGND VGND VPWR VPWR _4548_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7266_ _7265_/A _7265_/B _7265_/C VGND VGND VPWR VPWR _7377_/C sky130_fd_sc_hd__a21o_2
X_9005_ _8979_/A _8979_/B _8980_/A VGND VGND VPWR VPWR _9006_/A sky130_fd_sc_hd__o21ai_1
X_7197_ _7150_/A _7149_/A _7149_/B VGND VGND VPWR VPWR _7203_/A sky130_fd_sc_hd__o21ba_1
X_6217_ _6218_/A _6218_/B _6218_/C VGND VGND VPWR VPWR _6302_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6148_/A _6148_/B _6148_/C VGND VGND VPWR VPWR _6163_/C sky130_fd_sc_hd__nand3_1
XFILLER_57_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6079_ _9171_/Q VGND VGND VPWR VPWR _7453_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ _5450_/A VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5381_ _5367_/X _5653_/A _5377_/X _5379_/Y _5380_/X VGND VGND VPWR VPWR _5381_/X
+ sky130_fd_sc_hd__a221o_1
X_7120_ _7006_/A _7119_/C _7119_/D _7506_/B VGND VGND VPWR VPWR _7121_/B sky130_fd_sc_hd__a22oi_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7051_ _7076_/A _7076_/B VGND VGND VPWR VPWR _7053_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A VGND VGND VPWR VPWR _9208_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6002_ _6126_/B VGND VGND VPWR VPWR _9052_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7953_ _7952_/A _7952_/B _7952_/C VGND VGND VPWR VPWR _8029_/A sky130_fd_sc_hd__a21oi_2
X_6904_ _6781_/A _6780_/B _6780_/A VGND VGND VPWR VPWR _7033_/A sky130_fd_sc_hd__o21ba_1
X_7884_ _8587_/B VGND VGND VPWR VPWR _8780_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6835_ _6834_/A _6834_/B _6834_/C VGND VGND VPWR VPWR _6835_/X sky130_fd_sc_hd__a21o_1
X_6766_ _6766_/A _6766_/B VGND VGND VPWR VPWR _6767_/C sky130_fd_sc_hd__xnor2_1
X_8505_ _9004_/B VGND VGND VPWR VPWR _9025_/B sky130_fd_sc_hd__buf_4
X_5717_ _5712_/S _4541_/A _4889_/A VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__a21o_1
X_6697_ _6405_/B _7222_/C _7222_/D _6859_/A VGND VGND VPWR VPWR _6698_/B sky130_fd_sc_hd__a22o_1
X_8436_ _8664_/C VGND VGND VPWR VPWR _8844_/B sky130_fd_sc_hd__clkbuf_2
X_5648_ _5484_/A _5678_/A _5646_/X _5647_/Y _4541_/A VGND VGND VPWR VPWR _5648_/X
+ sky130_fd_sc_hd__a221o_1
X_8367_ _8379_/A _8450_/C _8450_/D _8452_/A VGND VGND VPWR VPWR _8370_/A sky130_fd_sc_hd__a22oi_1
X_5579_ _5509_/X _5577_/X _5674_/S VGND VGND VPWR VPWR _5579_/X sky130_fd_sc_hd__mux2_1
X_8298_ _8299_/A _8299_/B _8299_/C VGND VGND VPWR VPWR _8393_/B sky130_fd_sc_hd__o21a_1
X_7318_ _7449_/A _7449_/B VGND VGND VPWR VPWR _7319_/C sky130_fd_sc_hd__xnor2_1
X_7249_ _7324_/A _7249_/B VGND VGND VPWR VPWR _7377_/A sky130_fd_sc_hd__xnor2_2
XFILLER_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 A[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4950_ _4950_/A _4950_/B VGND VGND VPWR VPWR _4951_/B sky130_fd_sc_hd__nor2_1
X_4881_ _4608_/B _4838_/Y _4876_/Y _4877_/Y _5606_/A VGND VGND VPWR VPWR _4881_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6620_ _6618_/X _6619_/Y _6548_/C _6550_/A VGND VGND VPWR VPWR _6640_/B sky130_fd_sc_hd__a211o_1
X_6551_ _6551_/A _6551_/B VGND VGND VPWR VPWR _6643_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5502_ _5402_/X _5501_/X _5552_/S VGND VGND VPWR VPWR _5502_/X sky130_fd_sc_hd__mux2_1
X_6482_ _6483_/B _6483_/C _6483_/A VGND VGND VPWR VPWR _6646_/A sky130_fd_sc_hd__o21ai_2
X_8221_ _8221_/A _8221_/B VGND VGND VPWR VPWR _8223_/A sky130_fd_sc_hd__xor2_1
X_5433_ _5433_/A VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8152_ _8519_/A _8595_/A VGND VGND VPWR VPWR _8153_/B sky130_fd_sc_hd__nand2_1
X_5364_ _5364_/A VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7103_/A _7103_/B VGND VGND VPWR VPWR _7104_/C sky130_fd_sc_hd__nand2_1
X_8083_ _8083_/A _7995_/A VGND VGND VPWR VPWR _8100_/B sky130_fd_sc_hd__or2b_1
XFILLER_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5295_ _4599_/A _5485_/A _5378_/A VGND VGND VPWR VPWR _5295_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_87_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7034_ _7034_/A _6911_/B VGND VGND VPWR VPWR _7048_/B sky130_fd_sc_hd__or2b_1
XFILLER_67_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8985_ _8985_/A _8985_/B VGND VGND VPWR VPWR _8986_/B sky130_fd_sc_hd__or2_1
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7936_ _7848_/A _7850_/B _7848_/B VGND VGND VPWR VPWR _7942_/A sky130_fd_sc_hd__o21ba_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7867_ _8674_/A VGND VGND VPWR VPWR _8733_/A sky130_fd_sc_hd__buf_2
X_6818_ _7295_/C VGND VGND VPWR VPWR _7562_/A sky130_fd_sc_hd__clkbuf_2
X_7798_ _7689_/A _8639_/B _7690_/A _7688_/B VGND VGND VPWR VPWR _7911_/A sky130_fd_sc_hd__a31o_1
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6749_ _6747_/A _6952_/A _6748_/Y VGND VGND VPWR VPWR _6849_/A sky130_fd_sc_hd__o21ai_1
X_8419_ _8419_/A _8419_/B _8419_/C VGND VGND VPWR VPWR _8420_/B sky130_fd_sc_hd__nor3_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5080_ _5080_/A _5080_/B _5080_/C VGND VGND VPWR VPWR _5080_/X sky130_fd_sc_hd__or3_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8770_ _8770_/A _8770_/B VGND VGND VPWR VPWR _8771_/B sky130_fd_sc_hd__nor2_1
X_5982_ _5985_/D VGND VGND VPWR VPWR _6424_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7721_ _7801_/A VGND VGND VPWR VPWR _7724_/C sky130_fd_sc_hd__inv_2
X_4933_ _4933_/A _4937_/B VGND VGND VPWR VPWR _4933_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_13 _9133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7652_ _7651_/A _7651_/B _7651_/C VGND VGND VPWR VPWR _7772_/A sky130_fd_sc_hd__o21a_1
X_4864_ _4864_/A _4960_/A VGND VGND VPWR VPWR _5054_/S sky130_fd_sc_hd__nand2_2
XANTENNA_57 _9140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _7583_/A _7583_/B _7938_/C _7583_/D VGND VGND VPWR VPWR _7712_/A sky130_fd_sc_hd__and4_1
X_6603_ _6532_/A _6531_/A _6531_/B VGND VGND VPWR VPWR _6695_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_35 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _9198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _5571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4795_ _5733_/S _4960_/A _4794_/X VGND VGND VPWR VPWR _4795_/Y sky130_fd_sc_hd__o21ai_1
X_6534_ _7506_/A _7506_/B _7822_/B _6663_/C VGND VGND VPWR VPWR _6536_/A sky130_fd_sc_hd__and4_1
X_6465_ _6464_/A _6483_/C _6462_/Y _6551_/A VGND VGND VPWR VPWR _6465_/X sky130_fd_sc_hd__a2bb2o_1
X_8204_ _8203_/A _8203_/B _8203_/C VGND VGND VPWR VPWR _8318_/A sky130_fd_sc_hd__a21oi_2
X_5416_ _5266_/X _5122_/X _5413_/X _5415_/Y _4550_/A VGND VGND VPWR VPWR _5416_/X
+ sky130_fd_sc_hd__a221o_1
X_6396_ _7148_/D VGND VGND VPWR VPWR _7728_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_9184_ _9220_/CLK _9184_/D VGND VGND VPWR VPWR _9184_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8135_ _8135_/A _8135_/B VGND VGND VPWR VPWR _8211_/A sky130_fd_sc_hd__nand2_1
X_5347_ _5214_/X _5179_/X _5345_/X _5346_/Y _5001_/A VGND VGND VPWR VPWR _5347_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8066_ _8064_/X _8217_/A _7948_/B _7951_/B VGND VGND VPWR VPWR _8111_/A sky130_fd_sc_hd__o211a_1
X_5278_ _5656_/A VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__clkbuf_4
X_7017_ _7129_/A _7822_/B VGND VGND VPWR VPWR _7021_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8968_ _8920_/A _8920_/B _8921_/A VGND VGND VPWR VPWR _8968_/X sky130_fd_sc_hd__o21ba_1
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7919_ _7919_/A _7919_/B VGND VGND VPWR VPWR _8012_/A sky130_fd_sc_hd__xnor2_1
X_8899_ _8900_/A _8900_/B VGND VGND VPWR VPWR _8901_/A sky130_fd_sc_hd__or2_1
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput11 A[19] VGND VGND VPWR VPWR _9181_/D sky130_fd_sc_hd__clkbuf_1
X_4580_ _5559_/B VGND VGND VPWR VPWR _4580_/X sky130_fd_sc_hd__buf_2
Xinput22 A[29] VGND VGND VPWR VPWR _9191_/D sky130_fd_sc_hd__clkbuf_1
Xinput33 B[0] VGND VGND VPWR VPWR _9193_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 B[1] VGND VGND VPWR VPWR _9194_/D sky130_fd_sc_hd__clkbuf_1
Xinput55 B[2] VGND VGND VPWR VPWR _9195_/D sky130_fd_sc_hd__clkbuf_4
X_6250_ _6157_/B _6161_/B _6157_/A VGND VGND VPWR VPWR _6260_/A sky130_fd_sc_hd__o21ba_1
XFILLER_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6181_ _6268_/A _6181_/B VGND VGND VPWR VPWR _6264_/A sky130_fd_sc_hd__xnor2_1
X_5201_ _5743_/S VGND VGND VPWR VPWR _5365_/A sky130_fd_sc_hd__clkbuf_2
X_5132_ _5132_/A VGND VGND VPWR VPWR _5132_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5063_ _5059_/X _5060_/X _5062_/X _5164_/A VGND VGND VPWR VPWR _5063_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8822_ _8756_/A _9025_/B _8757_/A _8755_/B VGND VGND VPWR VPWR _8829_/B sky130_fd_sc_hd__a31oi_4
X_8753_ _8753_/A _8753_/B _8752_/Y VGND VGND VPWR VPWR _8755_/A sky130_fd_sc_hd__nor3b_1
X_5965_ _5965_/A _5965_/B _5965_/C VGND VGND VPWR VPWR _5968_/A sky130_fd_sc_hd__or3_1
X_8684_ _8684_/A _8684_/B VGND VGND VPWR VPWR _8686_/A sky130_fd_sc_hd__xor2_1
X_7704_ _7606_/A _7605_/A _7605_/B VGND VGND VPWR VPWR _7710_/A sky130_fd_sc_hd__o21ba_1
X_5896_ _5897_/A _5896_/B _9060_/A VGND VGND VPWR VPWR _5951_/B sky130_fd_sc_hd__or3b_1
X_4916_ _5054_/S _5052_/A _4915_/Y VGND VGND VPWR VPWR _4916_/X sky130_fd_sc_hd__a21o_1
X_7635_ _7635_/A _7635_/B VGND VGND VPWR VPWR _7740_/A sky130_fd_sc_hd__nand2_1
X_4847_ _4847_/A VGND VGND VPWR VPWR _4847_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7566_ _7569_/D VGND VGND VPWR VPWR _7566_/Y sky130_fd_sc_hd__clkinv_2
X_4778_ _4778_/A VGND VGND VPWR VPWR _5656_/B sky130_fd_sc_hd__buf_2
X_7497_ _7988_/B VGND VGND VPWR VPWR _8156_/C sky130_fd_sc_hd__clkbuf_2
X_6517_ _6257_/C _7148_/B _6424_/D _7148_/A VGND VGND VPWR VPWR _6518_/B sky130_fd_sc_hd__a22oi_1
X_6448_ _6894_/A _7006_/B _7327_/B _7152_/D VGND VGND VPWR VPWR _6451_/A sky130_fd_sc_hd__and4_1
X_9167_ _9210_/CLK _9167_/D VGND VGND VPWR VPWR _9167_/Q sky130_fd_sc_hd__dfxtp_2
X_6379_ _6473_/A _6379_/B VGND VGND VPWR VPWR _6480_/B sky130_fd_sc_hd__xor2_4
X_8118_ _8118_/A _8011_/A VGND VGND VPWR VPWR _8118_/X sky130_fd_sc_hd__or2b_1
XFILLER_102_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9098_ _9221_/CLK _9098_/D VGND VGND VPWR VPWR _9098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8049_ _8050_/B _8050_/C _8720_/A _8050_/A VGND VGND VPWR VPWR _8051_/A sky130_fd_sc_hd__a22oi_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5750_ _5402_/X _5484_/X _5749_/Y _4876_/A VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__o31a_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4701_/A _4828_/A VGND VGND VPWR VPWR _4705_/A sky130_fd_sc_hd__and2_2
X_5681_ _4783_/A _9089_/Q _4582_/A VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__a21o_1
X_7420_ _7421_/C _7696_/B _7418_/Y _7419_/X VGND VGND VPWR VPWR _7422_/A sky130_fd_sc_hd__o2bb2a_1
X_4632_ _5154_/A VGND VGND VPWR VPWR _5368_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7351_ _7351_/A _7351_/B VGND VGND VPWR VPWR _7352_/C sky130_fd_sc_hd__xnor2_1
X_4563_ _9096_/Q VGND VGND VPWR VPWR _5727_/S sky130_fd_sc_hd__inv_2
X_6302_ _6302_/A _6302_/B VGND VGND VPWR VPWR _6303_/B sky130_fd_sc_hd__nand2_1
X_7282_ _7403_/A _7282_/B VGND VGND VPWR VPWR _7284_/A sky130_fd_sc_hd__nor2_1
X_9021_ _8972_/A _8972_/B _8999_/A _8999_/B _9020_/Y VGND VGND VPWR VPWR _9022_/B
+ sky130_fd_sc_hd__o41a_1
X_6233_ _7307_/A VGND VGND VPWR VPWR _7146_/A sky130_fd_sc_hd__clkbuf_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6087_/A _6087_/B _6087_/C VGND VGND VPWR VPWR _6166_/C sky130_fd_sc_hd__a21bo_1
XFILLER_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6680_/B VGND VGND VPWR VPWR _7986_/A sky130_fd_sc_hd__clkbuf_4
X_5115_ _9089_/Q VGND VGND VPWR VPWR _5116_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5046_ _5067_/B _5046_/B VGND VGND VPWR VPWR _5046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8805_ _8805_/A _8731_/B VGND VGND VPWR VPWR _8806_/A sky130_fd_sc_hd__or2b_1
X_6997_ _9181_/Q VGND VGND VPWR VPWR _7259_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8736_ _8736_/A _8736_/B VGND VGND VPWR VPWR _8738_/A sky130_fd_sc_hd__xnor2_1
XFILLER_13_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5948_ _5948_/A _5948_/B _9064_/A VGND VGND VPWR VPWR _9062_/A sky130_fd_sc_hd__and3_1
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8667_ _8667_/A _8667_/B VGND VGND VPWR VPWR _8668_/C sky130_fd_sc_hd__xnor2_1
X_5879_ _7421_/C VGND VGND VPWR VPWR _7689_/A sky130_fd_sc_hd__clkbuf_2
X_7618_ _7472_/B _7618_/B VGND VGND VPWR VPWR _7618_/X sky130_fd_sc_hd__and2b_1
X_8598_ _8598_/A _8598_/B VGND VGND VPWR VPWR _8600_/A sky130_fd_sc_hd__xnor2_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7549_ _7549_/A _7549_/B VGND VGND VPWR VPWR _9090_/D sky130_fd_sc_hd__xnor2_1
X_9219_ _9219_/CLK _9219_/D VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6920_ _7569_/C _7849_/B VGND VGND VPWR VPWR _6924_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6851_ _6843_/A _6843_/B _6843_/C VGND VGND VPWR VPWR _6959_/A sky130_fd_sc_hd__a21bo_1
X_5802_ _7365_/A VGND VGND VPWR VPWR _7257_/A sky130_fd_sc_hd__buf_2
X_8521_ _8521_/A _8926_/B VGND VGND VPWR VPWR _8522_/B sky130_fd_sc_hd__nand2_1
X_6782_ _9178_/Q VGND VGND VPWR VPWR _7348_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5733_ _5214_/A _5732_/X _5733_/S VGND VGND VPWR VPWR _5733_/X sky130_fd_sc_hd__mux2_1
X_8452_ _8452_/A VGND VGND VPWR VPWR _8639_/A sky130_fd_sc_hd__clkbuf_2
X_5664_ _4650_/A _4716_/A _5662_/X _5663_/Y _4774_/A VGND VGND VPWR VPWR _5664_/X
+ sky130_fd_sc_hd__a221o_1
X_8383_ _8464_/B VGND VGND VPWR VPWR _8675_/A sky130_fd_sc_hd__clkbuf_2
X_5595_ _4573_/A _5385_/A _5175_/A VGND VGND VPWR VPWR _5595_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7403_ _7403_/A _7403_/B _7544_/A VGND VGND VPWR VPWR _7411_/A sky130_fd_sc_hd__and3_1
X_4615_ _5737_/S VGND VGND VPWR VPWR _5354_/S sky130_fd_sc_hd__buf_2
X_7334_ _7334_/A _7334_/B VGND VGND VPWR VPWR _7476_/B sky130_fd_sc_hd__xnor2_1
X_4546_ _9103_/Q VGND VGND VPWR VPWR _4721_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7265_ _7265_/A _7265_/B _7265_/C VGND VGND VPWR VPWR _7377_/B sky130_fd_sc_hd__nand3_1
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9004_ _9004_/A _9004_/B VGND VGND VPWR VPWR _9008_/A sky130_fd_sc_hd__nand2_1
X_7196_ _7421_/C _7940_/B _7085_/B _7084_/B VGND VGND VPWR VPWR _7204_/A sky130_fd_sc_hd__a31o_1
X_6216_ _6301_/A _6301_/B VGND VGND VPWR VPWR _6218_/C sky130_fd_sc_hd__xnor2_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6148_/A _6148_/B _6148_/C VGND VGND VPWR VPWR _6163_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6078_ _6256_/A VGND VGND VPWR VPWR _6500_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5029_ _9127_/Q _9119_/Q VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8719_ _8542_/B _8664_/D _8516_/B _8542_/A VGND VGND VPWR VPWR _8722_/A sky130_fd_sc_hd__a22oi_2
XFILLER_41_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5380_ _5382_/A VGND VGND VPWR VPWR _5380_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7050_ _7050_/A _7104_/A VGND VGND VPWR VPWR _7076_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6001_ _6047_/B _6001_/B VGND VGND VPWR VPWR _6126_/B sky130_fd_sc_hd__xor2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7952_ _7952_/A _7952_/B _7952_/C VGND VGND VPWR VPWR _7952_/X sky130_fd_sc_hd__and3_1
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6903_ _6802_/A _6801_/B _6801_/A VGND VGND VPWR VPWR _7034_/A sky130_fd_sc_hd__o21ba_1
XFILLER_54_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7883_ _8349_/B VGND VGND VPWR VPWR _8587_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6834_ _6834_/A _6834_/B _6834_/C VGND VGND VPWR VPWR _6836_/A sky130_fd_sc_hd__and3_1
X_6765_ _6917_/B _6765_/B VGND VGND VPWR VPWR _6766_/B sky130_fd_sc_hd__xnor2_1
X_8504_ _8504_/A _8504_/B VGND VGND VPWR VPWR _8513_/A sky130_fd_sc_hd__or2_1
X_5716_ _5676_/A _5714_/X _5715_/X VGND VGND VPWR VPWR _5716_/Y sky130_fd_sc_hd__a21oi_1
X_8435_ _8514_/A _8435_/B VGND VGND VPWR VPWR _8444_/A sky130_fd_sc_hd__xnor2_1
X_6696_ _6859_/A _7083_/A _7327_/C _7148_/D VGND VGND VPWR VPWR _6696_/X sky130_fd_sc_hd__and4_1
XFILLER_40_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5647_ _4870_/S _5271_/X _4883_/X VGND VGND VPWR VPWR _5647_/Y sky130_fd_sc_hd__a21oi_1
X_8366_ _8366_/A _8490_/A VGND VGND VPWR VPWR _8403_/A sky130_fd_sc_hd__nor2_1
X_5578_ _5697_/S VGND VGND VPWR VPWR _5674_/S sky130_fd_sc_hd__clkbuf_2
X_8297_ _8297_/A _8378_/B VGND VGND VPWR VPWR _8299_/C sky130_fd_sc_hd__xnor2_1
X_7317_ _7317_/A _7317_/B VGND VGND VPWR VPWR _7449_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7248_ _7248_/A _7340_/A VGND VGND VPWR VPWR _7249_/B sky130_fd_sc_hd__and2_1
XFILLER_49_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7179_ _7289_/A _7179_/B VGND VGND VPWR VPWR _7182_/B sky130_fd_sc_hd__and2_1
XFILLER_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 A[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4880_ _4880_/A VGND VGND VPWR VPWR _5606_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6550_ _6550_/A _6550_/B VGND VGND VPWR VPWR _6643_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5501_ _5364_/X _4769_/A _5499_/X _5500_/Y VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__a22o_1
X_6481_ _6481_/A _6481_/B VGND VGND VPWR VPWR _6557_/A sky130_fd_sc_hd__or2_1
X_8220_ _8220_/A _8816_/B VGND VGND VPWR VPWR _8221_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5432_ _5432_/A VGND VGND VPWR VPWR _5433_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8151_ _8151_/A _8151_/B VGND VGND VPWR VPWR _8153_/A sky130_fd_sc_hd__nor2_1
X_5363_ _5339_/X _5202_/X _5204_/X _5360_/X _5362_/X VGND VGND VPWR VPWR _9134_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7102_ _7102_/A _7102_/B _7215_/A VGND VGND VPWR VPWR _7103_/B sky130_fd_sc_hd__or3_2
X_8082_ _8082_/A _8082_/B VGND VGND VPWR VPWR _8105_/A sky130_fd_sc_hd__and2_1
XFILLER_99_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5294_ _5160_/A _5532_/A _5292_/X _5293_/Y _5410_/A VGND VGND VPWR VPWR _5294_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7033_ _7033_/A _6910_/B VGND VGND VPWR VPWR _7048_/A sky130_fd_sc_hd__or2b_1
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8984_ _8985_/A _8985_/B VGND VGND VPWR VPWR _9006_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7935_ _8177_/A _8185_/A _7935_/C VGND VGND VPWR VPWR _7944_/B sky130_fd_sc_hd__and3_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7866_ _8150_/D VGND VGND VPWR VPWR _8674_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6817_ _6817_/A _6817_/B VGND VGND VPWR VPWR _6834_/B sky130_fd_sc_hd__or2_1
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7797_ _7797_/A _7797_/B VGND VGND VPWR VPWR _9092_/D sky130_fd_sc_hd__xnor2_1
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6748_ _6748_/A _6748_/B VGND VGND VPWR VPWR _6748_/Y sky130_fd_sc_hd__nand2_1
X_6679_ _6679_/A VGND VGND VPWR VPWR _8038_/A sky130_fd_sc_hd__buf_2
X_8418_ _8418_/A VGND VGND VPWR VPWR _8420_/A sky130_fd_sc_hd__inv_2
X_8349_ _8349_/A _8349_/B _8349_/C VGND VGND VPWR VPWR _8349_/X sky130_fd_sc_hd__and3_1
XFILLER_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A VGND VGND VPWR VPWR _9116_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5981_ _9200_/Q VGND VGND VPWR VPWR _5985_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7720_ _7621_/C _7622_/B _7717_/X _7718_/Y VGND VGND VPWR VPWR _7801_/A sky130_fd_sc_hd__a211oi_2
XFILLER_52_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4932_ _4933_/A _4937_/B VGND VGND VPWR VPWR _4932_/X sky130_fd_sc_hd__or2_2
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7651_ _7651_/A _7651_/B _7651_/C VGND VGND VPWR VPWR _7653_/A sky130_fd_sc_hd__nor3_1
XANTENNA_14 _9133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6602_ _6601_/A _6601_/B _6601_/C VGND VGND VPWR VPWR _6691_/A sky130_fd_sc_hd__a21o_2
X_4863_ _4586_/A _4838_/Y _4859_/X _4862_/X VGND VGND VPWR VPWR _4863_/X sky130_fd_sc_hd__a211o_1
X_7582_ _7923_/B _8050_/C _8050_/D _6679_/A VGND VGND VPWR VPWR _7584_/A sky130_fd_sc_hd__a22oi_1
XANTENNA_36 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _9198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _5213_/A _4787_/B _4792_/X _4793_/Y _5071_/A VGND VGND VPWR VPWR _4794_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_25 _8780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _9140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _6593_/A _7728_/C VGND VGND VPWR VPWR _6537_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6464_ _6464_/A _6483_/C _6462_/Y _6551_/A VGND VGND VPWR VPWR _6551_/B sky130_fd_sc_hd__or4bb_1
X_8203_ _8203_/A _8203_/B _8203_/C VGND VGND VPWR VPWR _8203_/X sky130_fd_sc_hd__and3_1
X_5415_ _5382_/X _5189_/X _5414_/X VGND VGND VPWR VPWR _5415_/Y sky130_fd_sc_hd__a21oi_1
X_9183_ _9208_/CLK _9183_/D VGND VGND VPWR VPWR _9183_/Q sky130_fd_sc_hd__dfxtp_2
X_6395_ _9206_/Q VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__clkbuf_2
X_8134_ _8032_/A _9004_/B _8033_/A _8031_/B VGND VGND VPWR VPWR _8234_/A sky130_fd_sc_hd__a31o_1
X_5346_ _5003_/X _5131_/A _5135_/A VGND VGND VPWR VPWR _5346_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8065_ _8064_/A _8064_/B _8064_/C VGND VGND VPWR VPWR _8217_/A sky130_fd_sc_hd__a21oi_2
X_5277_ _9086_/Q VGND VGND VPWR VPWR _5656_/A sky130_fd_sc_hd__clkinv_2
XFILLER_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7016_ _7016_/A _7610_/C _7503_/C VGND VGND VPWR VPWR _7022_/A sky130_fd_sc_hd__and3_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8967_ _8967_/A VGND VGND VPWR VPWR _8967_/Y sky130_fd_sc_hd__inv_2
X_7918_ _7918_/A _8909_/B VGND VGND VPWR VPWR _7919_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8898_ _8949_/A _8898_/B VGND VGND VPWR VPWR _8900_/B sky130_fd_sc_hd__and2_1
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7849_ _8268_/A _7849_/B VGND VGND VPWR VPWR _7850_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 A[1] VGND VGND VPWR VPWR _9163_/D sky130_fd_sc_hd__clkbuf_1
Xinput45 B[20] VGND VGND VPWR VPWR _9213_/D sky130_fd_sc_hd__clkbuf_1
Xinput34 B[10] VGND VGND VPWR VPWR _9203_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 A[2] VGND VGND VPWR VPWR _9164_/D sky130_fd_sc_hd__buf_2
Xinput56 B[30] VGND VGND VPWR VPWR _9223_/D sky130_fd_sc_hd__clkbuf_1
X_5200_ _5200_/A VGND VGND VPWR VPWR _5200_/X sky130_fd_sc_hd__clkbuf_2
X_6180_ _6267_/A _6180_/B VGND VGND VPWR VPWR _6181_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5131_ _5131_/A VGND VGND VPWR VPWR _5581_/A sky130_fd_sc_hd__clkbuf_4
X_5062_ _4833_/A _5046_/Y _5061_/X _4598_/A VGND VGND VPWR VPWR _5062_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8821_ _8821_/A _8878_/A VGND VGND VPWR VPWR _8829_/A sky130_fd_sc_hd__or2_1
X_8752_ _8756_/A _8981_/B _8684_/A _8751_/X VGND VGND VPWR VPWR _8752_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7703_ _7703_/A _7703_/B VGND VGND VPWR VPWR _7718_/A sky130_fd_sc_hd__or2_1
XFILLER_52_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5964_ _6447_/A _9166_/Q _9167_/Q _6667_/A VGND VGND VPWR VPWR _5965_/C sky130_fd_sc_hd__a22oi_2
XFILLER_40_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8683_ _8756_/A _8850_/B VGND VGND VPWR VPWR _8684_/B sky130_fd_sc_hd__nand2_1
X_4915_ _4915_/A _5044_/A VGND VGND VPWR VPWR _4915_/Y sky130_fd_sc_hd__nor2_1
X_5895_ _9059_/A _9059_/B VGND VGND VPWR VPWR _9060_/A sky130_fd_sc_hd__and2_1
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7634_ _7635_/A _7635_/B VGND VGND VPWR VPWR _7636_/A sky130_fd_sc_hd__or2_1
X_4846_ _4846_/A VGND VGND VPWR VPWR _4847_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7565_ _6922_/B _7419_/C _7694_/D _7419_/B VGND VGND VPWR VPWR _7569_/D sky130_fd_sc_hd__a22o_1
X_6516_ _6680_/A _7307_/B _6760_/A _6680_/B VGND VGND VPWR VPWR _6611_/A sky130_fd_sc_hd__and4_1
X_4777_ _9093_/Q _5449_/A VGND VGND VPWR VPWR _4778_/A sky130_fd_sc_hd__nor2_1
X_7496_ _7496_/A _7496_/B VGND VGND VPWR VPWR _7514_/B sky130_fd_sc_hd__and2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6447_ _6447_/A VGND VGND VPWR VPWR _6894_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9166_ _9214_/CLK _9166_/D VGND VGND VPWR VPWR _9166_/Q sky130_fd_sc_hd__dfxtp_4
X_6378_ _6378_/A _6378_/B VGND VGND VPWR VPWR _6379_/B sky130_fd_sc_hd__nand2_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8117_ _8117_/A _8117_/B VGND VGND VPWR VPWR _8131_/A sky130_fd_sc_hd__or2_1
X_5329_ _4834_/A _5122_/X _5328_/X VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9097_ _9221_/CLK _9097_/D VGND VGND VPWR VPWR _9097_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8048_ _7960_/A _7963_/B _7960_/B VGND VGND VPWR VPWR _8054_/A sky130_fd_sc_hd__o21ba_1
XFILLER_75_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5680_ _9087_/Q _4579_/A _4658_/A _9086_/Q _5679_/Y VGND VGND VPWR VPWR _5680_/X
+ sky130_fd_sc_hd__o221a_1
X_4700_ _5187_/A VGND VGND VPWR VPWR _4769_/A sky130_fd_sc_hd__clkbuf_2
X_4631_ _5219_/A VGND VGND VPWR VPWR _5154_/A sky130_fd_sc_hd__buf_2
X_7350_ _7347_/Y _7490_/A _7349_/X VGND VGND VPWR VPWR _7351_/B sky130_fd_sc_hd__a21oi_1
X_4562_ _5729_/S VGND VGND VPWR VPWR _4870_/S sky130_fd_sc_hd__buf_2
X_6301_ _6301_/A _6301_/B VGND VGND VPWR VPWR _6302_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7281_ _7281_/A _7281_/B _7281_/C VGND VGND VPWR VPWR _7282_/B sky130_fd_sc_hd__nor3_1
X_9020_ _8964_/A _8999_/A _8999_/B VGND VGND VPWR VPWR _9020_/Y sky130_fd_sc_hd__o21bai_1
X_6232_ _6232_/A VGND VGND VPWR VPWR _7307_/A sky130_fd_sc_hd__buf_2
XFILLER_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6163_/A _6163_/B _6163_/C VGND VGND VPWR VPWR _6166_/B sky130_fd_sc_hd__nand3_1
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _7019_/B VGND VGND VPWR VPWR _6680_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5114_ _5114_/A _5114_/B VGND VGND VPWR VPWR _9159_/D sky130_fd_sc_hd__xnor2_4
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5072_/A VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__inv_2
XFILLER_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6996_ _7610_/C VGND VGND VPWR VPWR _7847_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8804_ _8804_/A _8804_/B VGND VGND VPWR VPWR _8863_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8735_ _8867_/A _8794_/B VGND VGND VPWR VPWR _8736_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5947_ _7645_/A _7531_/A _9067_/D VGND VGND VPWR VPWR _9064_/A sky130_fd_sc_hd__and3_1
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8666_ _8666_/A _8792_/A VGND VGND VPWR VPWR _8667_/B sky130_fd_sc_hd__nand2_1
X_7617_ _7616_/A _7616_/B _7616_/C VGND VGND VPWR VPWR _7621_/C sky130_fd_sc_hd__a21o_2
X_5878_ _7081_/A VGND VGND VPWR VPWR _7421_/C sky130_fd_sc_hd__clkbuf_2
X_8597_ _8597_/A _8597_/B VGND VGND VPWR VPWR _8598_/B sky130_fd_sc_hd__nand2_1
X_4829_ _4829_/A _4928_/A VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__or2_2
X_7548_ _7550_/B _7548_/B VGND VGND VPWR VPWR _7549_/B sky130_fd_sc_hd__nor2_1
X_7479_ _7485_/A VGND VGND VPWR VPWR _7873_/A sky130_fd_sc_hd__clkbuf_2
X_9218_ _9218_/CLK _9218_/D VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9149_ _9218_/CLK _9149_/D VGND VGND VPWR VPWR _9149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6850_ _6847_/A _6850_/B VGND VGND VPWR VPWR _6957_/A sky130_fd_sc_hd__nand2b_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5801_ _9194_/Q VGND VGND VPWR VPWR _7365_/A sky130_fd_sc_hd__buf_2
X_6781_ _6781_/A _6781_/B VGND VGND VPWR VPWR _6884_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8520_ _8520_/A _8520_/B VGND VGND VPWR VPWR _8523_/A sky130_fd_sc_hd__xnor2_1
X_5732_ _4789_/A _5731_/X _5732_/S VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__mux2_1
X_8451_ _8451_/A _8451_/B VGND VGND VPWR VPWR _8456_/A sky130_fd_sc_hd__nor2_1
X_5663_ _5558_/A _5214_/A _5000_/A VGND VGND VPWR VPWR _5663_/Y sky130_fd_sc_hd__a21oi_1
X_8382_ _8240_/A _8242_/B _8240_/B VGND VGND VPWR VPWR _8391_/A sky130_fd_sc_hd__o21ba_1
X_5594_ _5314_/A _5414_/A _5592_/X _5593_/Y _5173_/A VGND VGND VPWR VPWR _5594_/X
+ sky130_fd_sc_hd__a221o_1
X_7402_ _7403_/B _7544_/A _7403_/A VGND VGND VPWR VPWR _7404_/A sky130_fd_sc_hd__a21oi_1
X_4614_ _9106_/Q VGND VGND VPWR VPWR _5737_/S sky130_fd_sc_hd__inv_2
X_7333_ _7333_/A _7333_/B VGND VGND VPWR VPWR _7334_/B sky130_fd_sc_hd__nor2_1
X_4545_ _4545_/A VGND VGND VPWR VPWR _5632_/A sky130_fd_sc_hd__clkbuf_2
X_7264_ _7357_/A _7357_/B VGND VGND VPWR VPWR _7265_/C sky130_fd_sc_hd__xnor2_1
X_9003_ _9002_/A _9002_/B _9025_/A _9029_/A VGND VGND VPWR VPWR _9009_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6215_ _6304_/A _6215_/B VGND VGND VPWR VPWR _6301_/B sky130_fd_sc_hd__xnor2_1
X_7195_ _7195_/A _7195_/B VGND VGND VPWR VPWR _7321_/A sky130_fd_sc_hd__xor2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6068_/A _6068_/C _6068_/B VGND VGND VPWR VPWR _6148_/C sky130_fd_sc_hd__a21bo_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6077_ _6754_/B _6313_/B _7706_/A _6313_/A VGND VGND VPWR VPWR _6081_/A sky130_fd_sc_hd__a22oi_1
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5028_ _5028_/A _5028_/B VGND VGND VPWR VPWR _9157_/D sky130_fd_sc_hd__xor2_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6979_ _7077_/B _7079_/B VGND VGND VPWR VPWR _6980_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8718_ _8832_/A _8949_/A _8667_/A _8665_/B VGND VGND VPWR VPWR _8728_/B sky130_fd_sc_hd__a31o_1
X_8649_ _8649_/A _8649_/B VGND VGND VPWR VPWR _8773_/A sky130_fd_sc_hd__xor2_1
XFILLER_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6000_ _6000_/A _6047_/A VGND VGND VPWR VPWR _6001_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7951_ _7951_/A _7951_/B VGND VGND VPWR VPWR _7952_/C sky130_fd_sc_hd__nand2_1
X_7882_ _8516_/B VGND VGND VPWR VPWR _8831_/B sky130_fd_sc_hd__buf_2
X_6902_ _6901_/A _6901_/B _6901_/C VGND VGND VPWR VPWR _7029_/A sky130_fd_sc_hd__a21o_2
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6833_ _6882_/B _6833_/B VGND VGND VPWR VPWR _6834_/C sky130_fd_sc_hd__xnor2_2
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6764_ _6704_/B _6706_/B _6704_/A VGND VGND VPWR VPWR _6765_/B sky130_fd_sc_hd__o21ba_1
X_8503_ _8419_/B _8420_/B _8500_/Y _8572_/A VGND VGND VPWR VPWR _8504_/B sky130_fd_sc_hd__o211a_1
X_6695_ _6695_/A _6609_/B VGND VGND VPWR VPWR _6710_/A sky130_fd_sc_hd__or2b_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5715_ _5557_/A _5678_/A _4541_/A VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a21o_1
X_8434_ _8521_/A _8844_/D _8351_/D _8349_/X VGND VGND VPWR VPWR _8435_/B sky130_fd_sc_hd__a31o_1
X_5646_ _5433_/A _4880_/A _5644_/X _5645_/Y _5271_/X VGND VGND VPWR VPWR _5646_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8365_ _8365_/A _8365_/B VGND VGND VPWR VPWR _8490_/A sky130_fd_sc_hd__nor2_1
X_5577_ _5484_/X _5575_/X _5673_/S VGND VGND VPWR VPWR _5577_/X sky130_fd_sc_hd__mux2_1
X_8296_ _8296_/A _8296_/B VGND VGND VPWR VPWR _8378_/B sky130_fd_sc_hd__xnor2_1
X_7316_ _7316_/A _7316_/B VGND VGND VPWR VPWR _7317_/B sky130_fd_sc_hd__or2_1
X_7247_ _7246_/A _7246_/B _7246_/C VGND VGND VPWR VPWR _7340_/A sky130_fd_sc_hd__o21ai_2
XFILLER_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7178_ _7177_/B _7287_/B _7177_/A VGND VGND VPWR VPWR _7179_/B sky130_fd_sc_hd__o21ai_1
XFILLER_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6129_ _6125_/A _6125_/B _6053_/B _6051_/B _6051_/A VGND VGND VPWR VPWR _6218_/A
+ sky130_fd_sc_hd__a2111o_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5500_ _4573_/X _5276_/X _4697_/A VGND VGND VPWR VPWR _5500_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6480_ _6480_/A _6480_/B _6560_/B VGND VGND VPWR VPWR _6480_/X sky130_fd_sc_hd__or3_1
X_5431_ _5402_/X _5365_/X _5366_/X _5429_/X _5430_/X VGND VGND VPWR VPWR _9136_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_99_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8150_ _8517_/A _8516_/A _8150_/C _8150_/D VGND VGND VPWR VPWR _8151_/B sky130_fd_sc_hd__and4_1
X_5362_ _5362_/A _5482_/B VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__or2_1
X_8081_ _8081_/A _8081_/B VGND VGND VPWR VPWR _8082_/B sky130_fd_sc_hd__or2_1
X_7101_ _7102_/B _7215_/A _7102_/A VGND VGND VPWR VPWR _7103_/A sky130_fd_sc_hd__o21ai_1
XFILLER_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7032_ _6933_/A _6933_/B _7031_/X VGND VGND VPWR VPWR _7076_/A sky130_fd_sc_hd__a21oi_2
X_5293_ _5249_/A _5166_/Y _5258_/A VGND VGND VPWR VPWR _5293_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8983_ _8983_/A VGND VGND VPWR VPWR _8985_/B sky130_fd_sc_hd__inv_2
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7934_ _7826_/A _7934_/B VGND VGND VPWR VPWR _7946_/A sky130_fd_sc_hd__and2b_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7865_ _7865_/A _7865_/B VGND VGND VPWR VPWR _7891_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7796_ _7796_/A _7796_/B VGND VGND VPWR VPWR _7797_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6816_ _6814_/C _6814_/Y _6812_/Y _6813_/X VGND VGND VPWR VPWR _6945_/C sky130_fd_sc_hd__o211ai_4
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6747_ _6747_/A _6952_/A VGND VGND VPWR VPWR _9083_/D sky130_fd_sc_hd__xor2_1
X_6678_ _6592_/A _6591_/A _6591_/B VGND VGND VPWR VPWR _6751_/A sky130_fd_sc_hd__o21ba_1
X_8417_ _8419_/A _8419_/B _8419_/C VGND VGND VPWR VPWR _8418_/A sky130_fd_sc_hd__o21ai_1
X_5629_ _5583_/X _5627_/X _5698_/S VGND VGND VPWR VPWR _5629_/X sky130_fd_sc_hd__mux2_1
X_8348_ _8351_/D VGND VGND VPWR VPWR _8348_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8279_ _8279_/A VGND VGND VPWR VPWR _8498_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5980_ _7131_/A VGND VGND VPWR VPWR _6257_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4931_ _5140_/A _4980_/B _5007_/B _4861_/A VGND VGND VPWR VPWR _4931_/X sky130_fd_sc_hd__a31o_1
X_7650_ _7770_/C _7648_/Y _7649_/X VGND VGND VPWR VPWR _7651_/C sky130_fd_sc_hd__o21a_1
X_4862_ _4862_/A VGND VGND VPWR VPWR _4862_/X sky130_fd_sc_hd__clkbuf_2
X_6601_ _6601_/A _6601_/B _6601_/C VGND VGND VPWR VPWR _6614_/B sky130_fd_sc_hd__nand3_1
XANTENNA_15 _9133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _7461_/A _7460_/A _7460_/B VGND VGND VPWR VPWR _7588_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_37 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _9198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _4830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4793_ _4716_/A _4760_/X _4774_/A VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__a21oi_1
X_6532_ _6532_/A _6532_/B VGND VGND VPWR VPWR _6585_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_59 _9130_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6463_ _6347_/C _6350_/B _6460_/X _6461_/Y VGND VGND VPWR VPWR _6551_/A sky130_fd_sc_hd__a211o_1
X_9182_ _9210_/CLK _9182_/D VGND VGND VPWR VPWR _9182_/Q sky130_fd_sc_hd__dfxtp_1
X_8202_ _8202_/A _8202_/B VGND VGND VPWR VPWR _8203_/C sky130_fd_sc_hd__nand2_1
X_5414_ _5414_/A VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__clkbuf_2
X_8133_ _8949_/B VGND VGND VPWR VPWR _9004_/B sky130_fd_sc_hd__clkbuf_4
X_6394_ _7189_/C _7959_/A _8084_/A _7096_/A VGND VGND VPWR VPWR _6399_/A sky130_fd_sc_hd__a22oi_2
XFILLER_99_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5345_ _5215_/X _5172_/A _5343_/X _5344_/Y _5222_/X VGND VGND VPWR VPWR _5345_/X
+ sky130_fd_sc_hd__a221o_1
X_8064_ _8064_/A _8064_/B _8064_/C VGND VGND VPWR VPWR _8064_/X sky130_fd_sc_hd__and3_1
X_5276_ _5391_/A VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7015_ _6909_/A _6908_/A _6908_/B VGND VGND VPWR VPWR _7145_/A sky130_fd_sc_hd__o21ba_1
XFILLER_68_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8966_ _8966_/A _8966_/B VGND VGND VPWR VPWR _8967_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7917_ _7917_/A _7917_/B VGND VGND VPWR VPWR _7919_/A sky130_fd_sc_hd__nor2_1
X_8897_ _8897_/A _8944_/A VGND VGND VPWR VPWR _8900_/A sky130_fd_sc_hd__xnor2_1
X_7848_ _7848_/A _7848_/B VGND VGND VPWR VPWR _7850_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7779_ _7779_/A _7779_/B VGND VGND VPWR VPWR _7782_/A sky130_fd_sc_hd__xnor2_4
XFILLER_51_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 A[20] VGND VGND VPWR VPWR _9182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput35 B[11] VGND VGND VPWR VPWR _9204_/D sky130_fd_sc_hd__clkbuf_1
Xinput24 A[30] VGND VGND VPWR VPWR _9192_/D sky130_fd_sc_hd__clkbuf_1
Xinput46 B[21] VGND VGND VPWR VPWR _9214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput57 B[31] VGND VGND VPWR VPWR _9065_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5130_ _9080_/Q VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__buf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5061_ _4925_/A _4950_/B _5067_/A _5067_/B VGND VGND VPWR VPWR _5061_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8820_ _8819_/A _8819_/B _8819_/C VGND VGND VPWR VPWR _8878_/A sky130_fd_sc_hd__o21a_1
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8751_ _8682_/B _8751_/B VGND VGND VPWR VPWR _8751_/X sky130_fd_sc_hd__and2b_1
X_5963_ _9194_/Q _6232_/A VGND VGND VPWR VPWR _5965_/B sky130_fd_sc_hd__nand2_1
X_7702_ _7702_/A _7702_/B VGND VGND VPWR VPWR _7703_/B sky130_fd_sc_hd__and2_1
X_4914_ _4914_/A _4943_/B VGND VGND VPWR VPWR _5052_/A sky130_fd_sc_hd__nor2_2
X_8682_ _8751_/B _8682_/B VGND VGND VPWR VPWR _8684_/A sky130_fd_sc_hd__xnor2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5894_ _5948_/A VGND VGND VPWR VPWR _9059_/B sky130_fd_sc_hd__inv_2
X_7633_ _7633_/A _7633_/B VGND VGND VPWR VPWR _7635_/B sky130_fd_sc_hd__xnor2_1
X_4845_ _4845_/A _4845_/B VGND VGND VPWR VPWR _4845_/Y sky130_fd_sc_hd__nand2_2
X_7564_ _7443_/A _7443_/B _7446_/B VGND VGND VPWR VPWR _7684_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4776_ _4776_/A VGND VGND VPWR VPWR _5449_/A sky130_fd_sc_hd__inv_2
X_6515_ _7146_/A VGND VGND VPWR VPWR _7810_/C sky130_fd_sc_hd__buf_2
X_7495_ _7371_/B _7495_/B VGND VGND VPWR VPWR _7514_/A sky130_fd_sc_hd__and2b_1
X_6446_ _6593_/A _7938_/B VGND VGND VPWR VPWR _6452_/A sky130_fd_sc_hd__nand2_1
X_9165_ _9224_/CLK _9165_/D VGND VGND VPWR VPWR _9165_/Q sky130_fd_sc_hd__dfxtp_2
X_6377_ _6377_/A _6377_/B VGND VGND VPWR VPWR _6473_/A sky130_fd_sc_hd__xnor2_4
XFILLER_88_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8116_ _8116_/A _8116_/B VGND VGND VPWR VPWR _8117_/B sky130_fd_sc_hd__nor2_1
X_9096_ _9221_/CLK _9096_/D VGND VGND VPWR VPWR _9096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5328_ _4878_/A _5208_/X _5326_/X _5327_/Y _9105_/Q VGND VGND VPWR VPWR _5328_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8047_ _8279_/A _8467_/A _8047_/C VGND VGND VPWR VPWR _8056_/B sky130_fd_sc_hd__and3_1
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A VGND VGND VPWR VPWR _9222_/CLK sky130_fd_sc_hd__clkbuf_2
X_5259_ _5249_/X _5404_/A _5257_/Y _5258_/X VGND VGND VPWR VPWR _5259_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8949_ _8949_/A _8949_/B VGND VGND VPWR VPWR _8951_/B sky130_fd_sc_hd__and2_1
XFILLER_71_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _9096_/Q VGND VGND VPWR VPWR _5219_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6300_ _6300_/A _6300_/B VGND VGND VPWR VPWR _6303_/A sky130_fd_sc_hd__or2_1
X_4561_ _9098_/Q VGND VGND VPWR VPWR _5729_/S sky130_fd_sc_hd__inv_2
X_7280_ _7281_/B _7281_/C _7281_/A VGND VGND VPWR VPWR _7403_/A sky130_fd_sc_hd__o21a_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6231_ _6231_/A _6329_/B _6231_/C VGND VGND VPWR VPWR _6332_/A sky130_fd_sc_hd__nand3_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6163_/B _6163_/C _6163_/A VGND VGND VPWR VPWR _6166_/A sky130_fd_sc_hd__a21o_1
XFILLER_69_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A _5113_/B VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__xnor2_2
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7293_/A _6859_/B _6257_/C _6424_/D VGND VGND VPWR VPWR _6097_/A sky130_fd_sc_hd__and4_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5044_ _5044_/A _5052_/B VGND VGND VPWR VPWR _5072_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8803_ _8803_/A _8803_/B VGND VGND VPWR VPWR _8804_/B sky130_fd_sc_hd__or2_1
X_6995_ _7346_/B VGND VGND VPWR VPWR _7610_/C sky130_fd_sc_hd__clkbuf_2
X_8734_ _8734_/A _8734_/B VGND VGND VPWR VPWR _8736_/A sky130_fd_sc_hd__nor2_1
X_5946_ _5946_/A VGND VGND VPWR VPWR _9067_/D sky130_fd_sc_hd__clkbuf_2
X_8665_ _8665_/A _8665_/B VGND VGND VPWR VPWR _8667_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5877_ _6974_/A VGND VGND VPWR VPWR _7081_/A sky130_fd_sc_hd__clkbuf_2
X_7616_ _7616_/A _7616_/B _7616_/C VGND VGND VPWR VPWR _7621_/B sky130_fd_sc_hd__nand3_1
X_4828_ _4828_/A _4828_/B _4828_/C VGND VGND VPWR VPWR _4939_/A sky130_fd_sc_hd__and3_1
X_8596_ _8596_/A _8596_/B VGND VGND VPWR VPWR _8598_/A sky130_fd_sc_hd__nor2_1
X_7547_ _7405_/A _7547_/B VGND VGND VPWR VPWR _7550_/B sky130_fd_sc_hd__and2b_1
X_4759_ _4759_/A _4824_/A VGND VGND VPWR VPWR _4866_/A sky130_fd_sc_hd__nor2_1
X_7478_ _7476_/X _7339_/B _7474_/Y _7475_/X VGND VGND VPWR VPWR _7522_/B sky130_fd_sc_hd__o211ai_4
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9217_ _9222_/CLK _9217_/D VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
X_6429_ _7696_/C _7485_/A VGND VGND VPWR VPWR _6430_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9148_ _9199_/CLK _9148_/D VGND VGND VPWR VPWR _9148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9079_ _9214_/CLK _9079_/D VGND VGND VPWR VPWR _9079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6780_ _6780_/A _6780_/B VGND VGND VPWR VPWR _6781_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5800_ _6014_/A VGND VGND VPWR VPWR _7293_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5731_ _5730_/X _9097_/Q _9100_/Q VGND VGND VPWR VPWR _5731_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8450_ _8527_/A _8597_/A _8450_/C _8450_/D VGND VGND VPWR VPWR _8451_/B sky130_fd_sc_hd__and4_1
X_5662_ _5286_/A _5222_/A _5660_/X _5661_/Y _5214_/A VGND VGND VPWR VPWR _5662_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8381_ _8527_/A _8832_/A _8296_/A _8294_/B VGND VGND VPWR VPWR _8392_/A sky130_fd_sc_hd__a31o_1
X_5593_ _5450_/A _5382_/A _4641_/A VGND VGND VPWR VPWR _5593_/Y sky130_fd_sc_hd__a21oi_1
X_4613_ _5754_/A _4876_/A _4602_/Y _4608_/X _5713_/S VGND VGND VPWR VPWR _4613_/X
+ sky130_fd_sc_hd__o221a_1
X_7401_ _7284_/C _7285_/B _7398_/Y _7399_/X VGND VGND VPWR VPWR _7544_/A sky130_fd_sc_hd__a211o_1
X_7332_ _9202_/Q _9203_/Q _9174_/Q _9175_/Q VGND VGND VPWR VPWR _7333_/B sky130_fd_sc_hd__and4_1
X_4544_ _5271_/A VGND VGND VPWR VPWR _4545_/A sky130_fd_sc_hd__clkbuf_2
X_7263_ _7263_/A _7356_/A VGND VGND VPWR VPWR _7357_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9002_ _9002_/A _9002_/B _9025_/A _9029_/A VGND VGND VPWR VPWR _9009_/A sky130_fd_sc_hd__or4bb_1
X_6214_ _6221_/A _6221_/B _6213_/Y VGND VGND VPWR VPWR _6215_/B sky130_fd_sc_hd__o21a_1
X_7194_ _7194_/A _8044_/B VGND VGND VPWR VPWR _7195_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6145_/A _6145_/B _6145_/C VGND VGND VPWR VPWR _6148_/B sky130_fd_sc_hd__nand3_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _7359_/A VGND VGND VPWR VPWR _6313_/A sky130_fd_sc_hd__clkbuf_2
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5027_ _5510_/A _4915_/A _4971_/B _5026_/X _5506_/A VGND VGND VPWR VPWR _5028_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_72_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8717_ _8717_/A VGND VGND VPWR VPWR _8949_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _7295_/C _7309_/B _6978_/C VGND VGND VPWR VPWR _7079_/B sky130_fd_sc_hd__and3_1
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5929_ _5930_/A _5930_/B _5930_/C VGND VGND VPWR VPWR _5929_/X sky130_fd_sc_hd__a21o_1
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8648_ _8648_/A _8648_/B VGND VGND VPWR VPWR _8649_/B sky130_fd_sc_hd__nand2_1
X_8579_ _8579_/A _8578_/X VGND VGND VPWR VPWR _8582_/A sky130_fd_sc_hd__or2b_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7950_ _7950_/A _7950_/B VGND VGND VPWR VPWR _7951_/B sky130_fd_sc_hd__or2_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7881_ _8720_/B VGND VGND VPWR VPWR _8516_/B sky130_fd_sc_hd__clkbuf_2
X_6901_ _6901_/A _6901_/B _6901_/C VGND VGND VPWR VPWR _6913_/B sky130_fd_sc_hd__nand3_1
X_6832_ _6832_/A _6853_/A VGND VGND VPWR VPWR _6833_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6763_ _6763_/A _6763_/B VGND VGND VPWR VPWR _6917_/B sky130_fd_sc_hd__xnor2_2
X_8502_ _8500_/Y _8572_/A _8419_/B _8420_/B VGND VGND VPWR VPWR _8504_/A sky130_fd_sc_hd__a211oi_1
X_5714_ _5534_/A _5713_/X _5714_/S VGND VGND VPWR VPWR _5714_/X sky130_fd_sc_hd__mux2_1
X_6694_ _6579_/A _6579_/B _6693_/X VGND VGND VPWR VPWR _6817_/A sky130_fd_sc_hd__a21oi_2
X_8433_ _8521_/A _8926_/B _8522_/A _8432_/Y VGND VGND VPWR VPWR _8514_/A sky130_fd_sc_hd__a31o_1
X_5645_ _4566_/X _5385_/X _4880_/A VGND VGND VPWR VPWR _5645_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8364_ _8365_/A _8365_/B VGND VGND VPWR VPWR _8366_/A sky130_fd_sc_hd__and2_1
X_5576_ _5740_/S VGND VGND VPWR VPWR _5673_/S sky130_fd_sc_hd__clkbuf_2
X_8295_ _8379_/A _8782_/A VGND VGND VPWR VPWR _8296_/B sky130_fd_sc_hd__nand2_1
X_7315_ _7316_/A _7316_/B VGND VGND VPWR VPWR _7317_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7246_ _7246_/A _7246_/B _7246_/C VGND VGND VPWR VPWR _7248_/A sky130_fd_sc_hd__or3_1
X_7177_ _7177_/A _7177_/B _7287_/B VGND VGND VPWR VPWR _7289_/A sky130_fd_sc_hd__or3_2
X_6128_ _6128_/A _6128_/B VGND VGND VPWR VPWR _9076_/D sky130_fd_sc_hd__xnor2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6702_/B VGND VGND VPWR VPWR _7148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5430_ _5430_/A _5482_/B VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__or2_1
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5361_ _5506_/A VGND VGND VPWR VPWR _5482_/B sky130_fd_sc_hd__clkbuf_1
X_8080_ _8081_/A _8081_/B VGND VGND VPWR VPWR _8082_/A sky130_fd_sc_hd__nand2_1
X_5292_ _4862_/X _5482_/A _5290_/X _5291_/Y _4841_/A VGND VGND VPWR VPWR _5292_/X
+ sky130_fd_sc_hd__a221o_1
X_7100_ _7281_/A _7100_/B VGND VGND VPWR VPWR _7102_/A sky130_fd_sc_hd__or2_1
X_7031_ _6932_/B _7031_/B VGND VGND VPWR VPWR _7031_/X sky130_fd_sc_hd__and2b_1
XFILLER_67_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8982_ _8982_/A _8982_/B VGND VGND VPWR VPWR _8983_/A sky130_fd_sc_hd__xnor2_1
X_7933_ _7933_/A _7933_/B VGND VGND VPWR VPWR _7950_/A sky130_fd_sc_hd__or2_1
XFILLER_67_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7864_ _7920_/A _7920_/B VGND VGND VPWR VPWR _7894_/A sky130_fd_sc_hd__xnor2_2
XFILLER_82_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6815_ _6812_/Y _6813_/X _6814_/C _6814_/Y VGND VGND VPWR VPWR _6945_/B sky130_fd_sc_hd__a211o_1
X_7795_ _7795_/A _7795_/B _7795_/C VGND VGND VPWR VPWR _7796_/A sky130_fd_sc_hd__and3_1
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6746_ _6748_/A _6748_/B VGND VGND VPWR VPWR _6952_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6677_ _6606_/B _6608_/B _6606_/A VGND VGND VPWR VPWR _6752_/A sky130_fd_sc_hd__o21ba_1
X_8416_ _8416_/A _8416_/B VGND VGND VPWR VPWR _8419_/C sky130_fd_sc_hd__xor2_1
X_5628_ _5628_/A VGND VGND VPWR VPWR _5698_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_105_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8347_ _8156_/A _7769_/A _8349_/C VGND VGND VPWR VPWR _8351_/D sky130_fd_sc_hd__a21o_1
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5559_ _9082_/Q _5559_/B VGND VGND VPWR VPWR _5559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8278_ _8278_/A _8278_/B VGND VGND VPWR VPWR _8282_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7229_ _7342_/A _7342_/B VGND VGND VPWR VPWR _7231_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4930_ _4930_/A VGND VGND VPWR VPWR _5007_/B sky130_fd_sc_hd__inv_2
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4861_ _4861_/A VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6600_ _6659_/A _6659_/B VGND VGND VPWR VPWR _6601_/C sky130_fd_sc_hd__xnor2_1
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 _9134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7580_ _8032_/A _8467_/A _7438_/A _7436_/B VGND VGND VPWR VPWR _7589_/A sky130_fd_sc_hd__a31o_1
XANTENNA_38 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 _5630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4792_ _4597_/A _4773_/Y _4788_/X _4791_/Y _4716_/A VGND VGND VPWR VPWR _4792_/X
+ sky130_fd_sc_hd__a221o_1
X_6531_ _6531_/A _6531_/B VGND VGND VPWR VPWR _6532_/B sky130_fd_sc_hd__nor2_1
XANTENNA_49 _9198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6462_ _6460_/X _6461_/Y _6347_/C _6350_/B VGND VGND VPWR VPWR _6462_/Y sky130_fd_sc_hd__o211ai_1
X_9181_ _9210_/CLK _9181_/D VGND VGND VPWR VPWR _9181_/Q sky130_fd_sc_hd__dfxtp_1
X_8201_ _8201_/A _8201_/B VGND VGND VPWR VPWR _8202_/B sky130_fd_sc_hd__or2_1
X_6393_ _7847_/C VGND VGND VPWR VPWR _8084_/A sky130_fd_sc_hd__clkbuf_4
X_5413_ _5367_/X _5124_/X _5411_/X _5412_/Y _5380_/X VGND VGND VPWR VPWR _5413_/X
+ sky130_fd_sc_hd__a221o_1
X_8132_ _8132_/A _8132_/B VGND VGND VPWR VPWR _8229_/B sky130_fd_sc_hd__nand2_1
X_5344_ _4862_/A _5248_/A _4591_/A VGND VGND VPWR VPWR _5344_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8063_ _8063_/A _8063_/B VGND VGND VPWR VPWR _8064_/C sky130_fd_sc_hd__nand2_1
X_5275_ _4883_/X _5208_/X _5270_/Y _5274_/Y _5020_/X VGND VGND VPWR VPWR _5275_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7014_ _7013_/A _7013_/B _7013_/C VGND VGND VPWR VPWR _7141_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8965_ _8965_/A VGND VGND VPWR VPWR _8966_/B sky130_fd_sc_hd__inv_2
XFILLER_83_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8896_ _8845_/A _8847_/B _8845_/B VGND VGND VPWR VPWR _8944_/A sky130_fd_sc_hd__o21ba_1
X_7916_ _7915_/A _7915_/B _7914_/Y VGND VGND VPWR VPWR _7917_/B sky130_fd_sc_hd__o21ba_1
X_7847_ _7847_/A _8050_/B _7847_/C _7847_/D VGND VGND VPWR VPWR _7848_/B sky130_fd_sc_hd__and4_1
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7778_ _7895_/A _7895_/B VGND VGND VPWR VPWR _7779_/B sky130_fd_sc_hd__xor2_4
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6729_ _7299_/A _8721_/A _8607_/B _6358_/A VGND VGND VPWR VPWR _6730_/C sky130_fd_sc_hd__a22o_1
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 A[21] VGND VGND VPWR VPWR _9183_/D sky130_fd_sc_hd__clkbuf_1
Xinput36 B[12] VGND VGND VPWR VPWR _9205_/D sky130_fd_sc_hd__clkbuf_2
Xinput25 A[31] VGND VGND VPWR VPWR _9065_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput58 B[3] VGND VGND VPWR VPWR _9196_/D sky130_fd_sc_hd__clkbuf_1
Xinput47 B[22] VGND VGND VPWR VPWR _9215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5060_ _4870_/S _5053_/Y _4872_/S VGND VGND VPWR VPWR _5060_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8750_ _8750_/A _8777_/B VGND VGND VPWR VPWR _8759_/A sky130_fd_sc_hd__xnor2_1
X_5962_ _9196_/Q _6667_/A _9166_/Q _9167_/Q VGND VGND VPWR VPWR _5965_/A sky130_fd_sc_hd__and4_1
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7701_ _7702_/A _7702_/B VGND VGND VPWR VPWR _7703_/A sky130_fd_sc_hd__nor2_1
X_4913_ _4913_/A _4913_/B VGND VGND VPWR VPWR _4943_/B sky130_fd_sc_hd__xnor2_2
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8681_ _8596_/A _8598_/B _8596_/B VGND VGND VPWR VPWR _8682_/B sky130_fd_sc_hd__o21ba_1
X_5893_ _5987_/A _5939_/B VGND VGND VPWR VPWR _5948_/A sky130_fd_sc_hd__or2_1
XFILLER_21_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7632_ _7873_/A _7748_/A VGND VGND VPWR VPWR _7633_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ _4845_/A _4950_/A VGND VGND VPWR VPWR _4844_/X sky130_fd_sc_hd__or2_2
X_7563_ _7563_/A _7563_/B VGND VGND VPWR VPWR _7683_/A sky130_fd_sc_hd__xor2_1
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4775_ _5728_/S VGND VGND VPWR VPWR _5621_/A sky130_fd_sc_hd__clkbuf_2
X_6514_ _6445_/A _6444_/A _6444_/B VGND VGND VPWR VPWR _6565_/A sky130_fd_sc_hd__o21ba_1
X_7494_ _7601_/A _7601_/B VGND VGND VPWR VPWR _7516_/A sky130_fd_sc_hd__xnor2_1
X_6445_ _6445_/A _6445_/B VGND VGND VPWR VPWR _6456_/A sky130_fd_sc_hd__xnor2_2
X_6376_ _6376_/A _6376_/B VGND VGND VPWR VPWR _6377_/B sky130_fd_sc_hd__nor2_2
X_9164_ _9220_/CLK _9164_/D VGND VGND VPWR VPWR _9164_/Q sky130_fd_sc_hd__dfxtp_1
X_8115_ _8116_/A _8116_/B VGND VGND VPWR VPWR _8117_/A sky130_fd_sc_hd__and2_1
X_5327_ _5173_/A _5273_/X _4878_/A VGND VGND VPWR VPWR _5327_/Y sky130_fd_sc_hd__a21oi_1
X_9095_ _9221_/CLK _9095_/D VGND VGND VPWR VPWR _9095_/Q sky130_fd_sc_hd__dfxtp_1
X_8046_ _7942_/A _8046_/B VGND VGND VPWR VPWR _8058_/A sky130_fd_sc_hd__and2b_1
X_5258_ _5258_/A VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5189_ _5634_/A VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__buf_4
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8948_ _8948_/A _8948_/B VGND VGND VPWR VPWR _8951_/A sky130_fd_sc_hd__and2_1
XFILLER_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8879_ _8921_/A _8879_/B VGND VGND VPWR VPWR _8966_/A sky130_fd_sc_hd__and2_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4560_ _4560_/A VGND VGND VPWR VPWR _5509_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6230_ _6231_/A _6329_/B _6231_/C VGND VGND VPWR VPWR _6245_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6161_/A _6161_/B VGND VGND VPWR VPWR _6163_/A sky130_fd_sc_hd__xnor2_4
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _9128_/Q _9120_/Q VGND VGND VPWR VPWR _5113_/B sky130_fd_sc_hd__xor2_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6092_ _6013_/A _6016_/B _6013_/B VGND VGND VPWR VPWR _6186_/A sky130_fd_sc_hd__o21ba_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A _5043_/B VGND VGND VPWR VPWR _5043_/Y sky130_fd_sc_hd__xnor2_1
X_8802_ _8803_/A _8803_/B VGND VGND VPWR VPWR _8804_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6994_ _6994_/A _6994_/B VGND VGND VPWR VPWR _7013_/B sky130_fd_sc_hd__nand2_1
X_8733_ _8733_/A _8792_/A _8842_/A _8733_/D VGND VGND VPWR VPWR _8734_/B sky130_fd_sc_hd__and4_1
X_5945_ _5945_/A _6358_/A VGND VGND VPWR VPWR _5946_/A sky130_fd_sc_hd__and2_1
X_8664_ _8664_/A _8664_/B _8664_/C _8664_/D VGND VGND VPWR VPWR _8665_/B sky130_fd_sc_hd__and4_1
X_5876_ _5881_/A _5892_/A VGND VGND VPWR VPWR _5885_/B sky130_fd_sc_hd__nand2_1
X_7615_ _7615_/A _7615_/B VGND VGND VPWR VPWR _7616_/C sky130_fd_sc_hd__xnor2_1
XFILLER_21_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _4943_/A _4827_/B VGND VGND VPWR VPWR _4856_/B sky130_fd_sc_hd__nand2_4
X_8595_ _8595_/A _8675_/A _8595_/C _8595_/D VGND VGND VPWR VPWR _8596_/B sky130_fd_sc_hd__and4_1
XFILLER_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7546_ _7553_/A _7553_/B VGND VGND VPWR VPWR _7549_/A sky130_fd_sc_hd__nor2_1
X_4758_ _4864_/A _4762_/A VGND VGND VPWR VPWR _4852_/A sky130_fd_sc_hd__nor2_2
X_7477_ _7474_/Y _7475_/X _7476_/X _7339_/B VGND VGND VPWR VPWR _7522_/A sky130_fd_sc_hd__a211o_1
X_4689_ _4691_/A _4864_/A VGND VGND VPWR VPWR _4701_/A sky130_fd_sc_hd__or2_1
X_6428_ _6607_/B VGND VGND VPWR VPWR _7485_/A sky130_fd_sc_hd__buf_2
X_9216_ _9216_/CLK _9216_/D VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_2
X_9147_ _9208_/CLK _9147_/D VGND VGND VPWR VPWR _9147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6359_ _6359_/A _7608_/A VGND VGND VPWR VPWR _6363_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9078_ _9214_/CLK _9078_/D VGND VGND VPWR VPWR _9078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8029_ _8029_/A _8029_/B _8028_/Y VGND VGND VPWR VPWR _8031_/A sky130_fd_sc_hd__nor3b_1
XFILLER_84_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5730_ _9096_/Q _5729_/X _5730_/S VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__mux2_1
X_5661_ _5424_/A _4839_/A _5222_/A VGND VGND VPWR VPWR _5661_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7400_ _7398_/Y _7399_/X _7284_/C _7285_/B VGND VGND VPWR VPWR _7403_/B sky130_fd_sc_hd__o211ai_1
X_8380_ _8724_/A VGND VGND VPWR VPWR _8832_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A VGND VGND VPWR VPWR _9219_/CLK sky130_fd_sc_hd__clkbuf_2
X_5592_ _5244_/A _5367_/A _5590_/X _5591_/Y _5132_/A VGND VGND VPWR VPWR _5592_/X
+ sky130_fd_sc_hd__a221o_1
X_4612_ _4966_/A VGND VGND VPWR VPWR _5713_/S sky130_fd_sc_hd__clkbuf_2
X_7331_ _7152_/C _7019_/C _9175_/Q _9202_/Q VGND VGND VPWR VPWR _7333_/A sky130_fd_sc_hd__a22oi_1
X_4543_ _5125_/A VGND VGND VPWR VPWR _5271_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7262_ _7122_/A _7121_/B _7121_/A VGND VGND VPWR VPWR _7356_/A sky130_fd_sc_hd__o21ba_1
X_9001_ _9001_/A _9001_/B VGND VGND VPWR VPWR _9108_/D sky130_fd_sc_hd__xnor2_1
X_6213_ _6213_/A _6213_/B VGND VGND VPWR VPWR _6213_/Y sky130_fd_sc_hd__nand2_1
X_7193_ _9214_/Q VGND VGND VPWR VPWR _8044_/B sky130_fd_sc_hd__buf_2
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6145_/B _6145_/C _6145_/A VGND VGND VPWR VPWR _6148_/A sky130_fd_sc_hd__a21o_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6075_ _7327_/A VGND VGND VPWR VPWR _7706_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _4687_/X _4980_/B _5024_/X _5025_/Y _4896_/A VGND VGND VPWR VPWR _5026_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6977_ _6700_/A _7824_/B _6978_/C VGND VGND VPWR VPWR _7077_/B sky130_fd_sc_hd__a21oi_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8716_ _8716_/A _9029_/B VGND VGND VPWR VPWR _8778_/A sky130_fd_sc_hd__nand2_1
X_5928_ _5961_/C _5928_/B VGND VGND VPWR VPWR _5930_/C sky130_fd_sc_hd__xnor2_2
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8647_ _8709_/A _8709_/B VGND VGND VPWR VPWR _8649_/A sky130_fd_sc_hd__xnor2_1
X_5859_ _5858_/A _5858_/B _5858_/C VGND VGND VPWR VPWR _5860_/B sky130_fd_sc_hd__a21o_1
X_8578_ _8575_/X _8648_/B _8504_/B _8513_/Y VGND VGND VPWR VPWR _8578_/X sky130_fd_sc_hd__a211o_1
X_7529_ _7526_/X _7665_/B _7528_/X _7386_/X VGND VGND VPWR VPWR _7538_/A sky130_fd_sc_hd__o211a_1
XFILLER_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7880_ _7880_/A _8349_/B VGND VGND VPWR VPWR _7997_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6900_ _6994_/A _6994_/B VGND VGND VPWR VPWR _6901_/C sky130_fd_sc_hd__xnor2_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6831_ _6831_/A _6831_/B VGND VGND VPWR VPWR _6832_/A sky130_fd_sc_hd__nor2_1
X_8501_ _8501_/A _8501_/B _8501_/C VGND VGND VPWR VPWR _8572_/A sky130_fd_sc_hd__or3_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6762_ _6762_/A _6762_/B VGND VGND VPWR VPWR _6763_/B sky130_fd_sc_hd__nor2_1
X_5713_ _4560_/A _5712_/X _5713_/S VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__mux2_1
X_6693_ _6578_/B _6693_/B VGND VGND VPWR VPWR _6693_/X sky130_fd_sc_hd__and2b_1
X_8432_ _8521_/A _8891_/B _8832_/B _6192_/X VGND VGND VPWR VPWR _8432_/Y sky130_fd_sc_hd__a22oi_1
X_5644_ _4587_/X _4643_/A _5642_/X _5643_/Y _5385_/X VGND VGND VPWR VPWR _5644_/X
+ sky130_fd_sc_hd__a221o_1
X_8363_ _8363_/A _8482_/B VGND VGND VPWR VPWR _8365_/B sky130_fd_sc_hd__xor2_1
X_7314_ _7204_/A _7204_/B _7313_/X VGND VGND VPWR VPWR _7316_/B sky130_fd_sc_hd__a21oi_1
X_5575_ _5461_/X _5574_/X _5575_/S VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8294_ _8294_/A _8294_/B VGND VGND VPWR VPWR _8296_/A sky130_fd_sc_hd__nor2_1
X_7245_ _7245_/A _7245_/B VGND VGND VPWR VPWR _7246_/C sky130_fd_sc_hd__xnor2_1
XFILLER_98_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7176_ _7176_/A _7176_/B _7287_/A VGND VGND VPWR VPWR _7287_/B sky130_fd_sc_hd__nor3_2
X_6127_ _6051_/B _6053_/B _6126_/X VGND VGND VPWR VPWR _6128_/B sky130_fd_sc_hd__o21ai_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6058_ _9169_/Q VGND VGND VPWR VPWR _6702_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5009_ _4861_/A _5054_/S _5052_/A _4839_/A VGND VGND VPWR VPWR _5009_/X sky130_fd_sc_hd__a31o_1
XFILLER_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5360_ _5315_/X _5358_/X _5481_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
X_5291_ _4586_/A _5370_/A _4862_/X VGND VGND VPWR VPWR _5291_/Y sky130_fd_sc_hd__a21oi_1
X_7030_ _7029_/A _7029_/B _7029_/C VGND VGND VPWR VPWR _7053_/C sky130_fd_sc_hd__a21oi_4
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8981_ _9004_/A _8981_/B VGND VGND VPWR VPWR _8982_/B sky130_fd_sc_hd__and2_1
XFILLER_82_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7932_ _7932_/A _7932_/B VGND VGND VPWR VPWR _7933_/B sky130_fd_sc_hd__and2_1
XFILLER_70_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7863_ _7863_/A _7952_/A VGND VGND VPWR VPWR _7920_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6814_ _6814_/A _6814_/B _6814_/C VGND VGND VPWR VPWR _6814_/Y sky130_fd_sc_hd__nor3_2
X_7794_ _7792_/Y _7794_/B VGND VGND VPWR VPWR _7797_/A sky130_fd_sc_hd__and2b_1
XFILLER_11_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6745_ _6750_/A _6745_/B VGND VGND VPWR VPWR _6748_/B sky130_fd_sc_hd__xnor2_1
X_8415_ _8415_/A _8639_/B VGND VGND VPWR VPWR _8416_/B sky130_fd_sc_hd__nand2_1
X_6676_ _6675_/A _6675_/B _6675_/C VGND VGND VPWR VPWR _6810_/A sky130_fd_sc_hd__a21o_2
X_5627_ _5754_/B _5626_/X _5674_/S VGND VGND VPWR VPWR _5627_/X sky130_fd_sc_hd__mux2_1
X_8346_ _8351_/C VGND VGND VPWR VPWR _8521_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5558_ _5558_/A VGND VGND VPWR VPWR _5558_/X sky130_fd_sc_hd__clkbuf_2
X_8277_ _8371_/A _8452_/A _8450_/C _8450_/D VGND VGND VPWR VPWR _8278_/B sky130_fd_sc_hd__and4_1
X_7228_ _7602_/A _7462_/A _7225_/Y _7335_/A VGND VGND VPWR VPWR _7342_/B sky130_fd_sc_hd__o2bb2a_1
X_5489_ _5368_/X _5210_/A _5487_/X _5488_/Y _5156_/X VGND VGND VPWR VPWR _5489_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_76_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7159_ _7159_/A _7159_/B VGND VGND VPWR VPWR _7160_/B sky130_fd_sc_hd__and2_1
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4860_ _9096_/Q VGND VGND VPWR VPWR _4861_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_17 _9134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _7359_/A _6530_/B _7822_/A _6886_/B VGND VGND VPWR VPWR _6531_/B sky130_fd_sc_hd__and4_1
XANTENNA_39 _9165_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _5581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4791_ _5058_/A _4960_/A _5214_/A VGND VGND VPWR VPWR _4791_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6461_ _6512_/B _6546_/A _6512_/A VGND VGND VPWR VPWR _6461_/Y sky130_fd_sc_hd__a21oi_1
X_8200_ _8201_/A _8201_/B VGND VGND VPWR VPWR _8202_/A sky130_fd_sc_hd__nand2_1
X_9180_ _9218_/CLK _9180_/D VGND VGND VPWR VPWR _9180_/Q sky130_fd_sc_hd__dfxtp_4
X_6392_ _7222_/D VGND VGND VPWR VPWR _7847_/C sky130_fd_sc_hd__clkbuf_2
X_5412_ _5247_/X _5184_/X _5378_/X VGND VGND VPWR VPWR _5412_/Y sky130_fd_sc_hd__a21oi_1
X_8131_ _8131_/A _8120_/B VGND VGND VPWR VPWR _8229_/A sky130_fd_sc_hd__or2b_1
X_5343_ _4585_/A _5166_/Y _5342_/X _5219_/X VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__a211o_1
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8062_ _8062_/A _8062_/B VGND VGND VPWR VPWR _8063_/B sky130_fd_sc_hd__or2_1
X_5274_ _5271_/X _5273_/X _4629_/A VGND VGND VPWR VPWR _5274_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7013_ _7013_/A _7013_/B _7013_/C VGND VGND VPWR VPWR _7027_/B sky130_fd_sc_hd__nand3_1
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8964_ _8964_/A _8963_/X VGND VGND VPWR VPWR _8972_/A sky130_fd_sc_hd__or2b_1
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8895_ _8895_/A _8895_/B VGND VGND VPWR VPWR _8897_/A sky130_fd_sc_hd__xnor2_1
X_7915_ _7915_/A _7915_/B _7914_/Y VGND VGND VPWR VPWR _7917_/A sky130_fd_sc_hd__nor3b_1
X_7846_ _8190_/A _7459_/D _8190_/B _7959_/A VGND VGND VPWR VPWR _7848_/A sky130_fd_sc_hd__a22oi_1
XFILLER_62_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7777_ _7657_/A _7657_/B _7776_/X VGND VGND VPWR VPWR _7895_/B sky130_fd_sc_hd__a21oi_4
X_4989_ _5032_/A _4989_/B VGND VGND VPWR VPWR _4991_/B sky130_fd_sc_hd__nand2_1
X_6728_ _8720_/A VGND VGND VPWR VPWR _8607_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6659_ _6659_/A _6659_/B VGND VGND VPWR VPWR _6675_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8329_ _8336_/A _8336_/B VGND VGND VPWR VPWR _8329_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 A[3] VGND VGND VPWR VPWR _9165_/D sky130_fd_sc_hd__clkbuf_4
Xinput15 A[22] VGND VGND VPWR VPWR _9184_/D sky130_fd_sc_hd__clkbuf_1
Xinput37 B[13] VGND VGND VPWR VPWR _9206_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 B[23] VGND VGND VPWR VPWR _9216_/D sky130_fd_sc_hd__clkbuf_1
Xinput59 B[4] VGND VGND VPWR VPWR _9197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5961_ _7194_/A _8071_/A _5961_/C VGND VGND VPWR VPWR _5997_/A sky130_fd_sc_hd__and3_1
X_8680_ _8680_/A _8680_/B VGND VGND VPWR VPWR _8751_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7700_ _7804_/A _9214_/Q VGND VGND VPWR VPWR _7702_/B sky130_fd_sc_hd__and2_1
X_4912_ _4957_/B VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__clkbuf_2
X_7631_ _7852_/C VGND VGND VPWR VPWR _7748_/A sky130_fd_sc_hd__clkbuf_2
X_5892_ _5892_/A _5892_/B VGND VGND VPWR VPWR _5939_/B sky130_fd_sc_hd__or2_1
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4843_ _4845_/B VGND VGND VPWR VPWR _4950_/A sky130_fd_sc_hd__clkbuf_2
X_7562_ _7562_/A _7804_/B VGND VGND VPWR VPWR _7563_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4774_ _4774_/A VGND VGND VPWR VPWR _5213_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7493_ _7600_/A _7493_/B VGND VGND VPWR VPWR _7601_/B sky130_fd_sc_hd__xnor2_1
X_6513_ _6425_/A _6430_/B _6425_/B VGND VGND VPWR VPWR _6566_/A sky130_fd_sc_hd__o21ba_1
X_6444_ _6444_/A _6444_/B VGND VGND VPWR VPWR _6445_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6375_ _6375_/A _6466_/A _6375_/C VGND VGND VPWR VPWR _6376_/B sky130_fd_sc_hd__and3_1
X_9163_ _9224_/CLK _9163_/D VGND VGND VPWR VPWR _9163_/Q sky130_fd_sc_hd__dfxtp_2
X_8114_ _8114_/A _8114_/B VGND VGND VPWR VPWR _8116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5326_ _5169_/A _5653_/A _5324_/X _5325_/Y _4548_/A VGND VGND VPWR VPWR _5326_/X
+ sky130_fd_sc_hd__a221o_1
X_9094_ _9221_/CLK _9094_/D VGND VGND VPWR VPWR _9094_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8045_ _8045_/A _8045_/B VGND VGND VPWR VPWR _8062_/A sky130_fd_sc_hd__xor2_1
X_5257_ _5154_/X _9075_/Q _5256_/X _5156_/X VGND VGND VPWR VPWR _5257_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_68_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5188_ _9085_/Q VGND VGND VPWR VPWR _5634_/A sky130_fd_sc_hd__clkinv_2
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8947_ _8947_/A _8947_/B VGND VGND VPWR VPWR _8948_/B sky130_fd_sc_hd__or2_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8878_ _8878_/A _8878_/B _8878_/C VGND VGND VPWR VPWR _8879_/B sky130_fd_sc_hd__or3_1
X_7829_ _7946_/B _7829_/B VGND VGND VPWR VPWR _7829_/X sky130_fd_sc_hd__or2_1
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _7309_/A _6775_/A VGND VGND VPWR VPWR _6161_/B sky130_fd_sc_hd__nand2_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _9126_/Q _9118_/Q _5032_/B _5035_/B _5031_/B VGND VGND VPWR VPWR _5113_/A
+ sky130_fd_sc_hd__a311oi_4
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6029_/B _6032_/B _6029_/A VGND VGND VPWR VPWR _6187_/A sky130_fd_sc_hd__o21ba_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _4915_/A _4971_/B _5028_/A VGND VGND VPWR VPWR _5043_/B sky130_fd_sc_hd__o21a_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8801_ _8801_/A _8865_/B VGND VGND VPWR VPWR _8803_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6993_ _6993_/A _6899_/A VGND VGND VPWR VPWR _7013_/A sky130_fd_sc_hd__or2b_1
XFILLER_53_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8732_ _8792_/A _8842_/A _8844_/C _8909_/A VGND VGND VPWR VPWR _8734_/A sky130_fd_sc_hd__a22oi_2
X_5944_ _7096_/A VGND VGND VPWR VPWR _6358_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8663_ _8831_/A _8841_/A _8351_/B _8780_/A VGND VGND VPWR VPWR _8665_/A sky130_fd_sc_hd__a22oi_1
XFILLER_61_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ _7647_/A _7509_/A _6858_/A _5922_/A VGND VGND VPWR VPWR _5892_/A sky130_fd_sc_hd__and4_2
X_7614_ _7742_/B _7614_/B VGND VGND VPWR VPWR _7615_/B sky130_fd_sc_hd__xnor2_1
X_8594_ _8675_/A _8792_/B _8792_/D _8538_/A VGND VGND VPWR VPWR _8596_/A sky130_fd_sc_hd__a22oi_1
X_4826_ _4836_/A _4845_/B VGND VGND VPWR VPWR _4827_/B sky130_fd_sc_hd__or2_1
XFILLER_21_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7545_ _7544_/A _7544_/B _7544_/C VGND VGND VPWR VPWR _7553_/B sky130_fd_sc_hd__a21oi_2
X_4757_ _4817_/S _4757_/B VGND VGND VPWR VPWR _4762_/A sky130_fd_sc_hd__nand2_1
X_7476_ _7336_/B _7476_/B VGND VGND VPWR VPWR _7476_/X sky130_fd_sc_hd__and2b_1
X_4688_ _4688_/A _4688_/B VGND VGND VPWR VPWR _4864_/A sky130_fd_sc_hd__nand2_1
X_6427_ _7419_/B VGND VGND VPWR VPWR _7696_/C sky130_fd_sc_hd__clkbuf_2
X_9215_ _9224_/CLK _9215_/D VGND VGND VPWR VPWR _9215_/Q sky130_fd_sc_hd__dfxtp_2
X_9146_ _9199_/CLK _9146_/D VGND VGND VPWR VPWR _9146_/Q sky130_fd_sc_hd__dfxtp_1
X_6358_ _6358_/A _8517_/A VGND VGND VPWR VPWR _6366_/A sky130_fd_sc_hd__nand2_1
X_5309_ _5200_/X _5307_/X _5428_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9077_ _9214_/CLK _9077_/D VGND VGND VPWR VPWR _9077_/Q sky130_fd_sc_hd__dfxtp_1
X_6289_ _6287_/Y _6288_/X _6207_/C _6210_/B VGND VGND VPWR VPWR _6292_/B sky130_fd_sc_hd__o211ai_1
XFILLER_75_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8028_ _7929_/A _7929_/B _7933_/B VGND VGND VPWR VPWR _8028_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5660_ _9090_/Q _5219_/A _5658_/X _5659_/Y _4839_/A VGND VGND VPWR VPWR _5660_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4611_ _5691_/S VGND VGND VPWR VPWR _4966_/A sky130_fd_sc_hd__clkbuf_2
X_5591_ _5394_/A _5410_/A _5378_/A VGND VGND VPWR VPWR _5591_/Y sky130_fd_sc_hd__a21oi_1
X_7330_ _7330_/A _9204_/Q VGND VGND VPWR VPWR _7334_/A sky130_fd_sc_hd__nand2_1
X_4542_ _9105_/Q VGND VGND VPWR VPWR _5125_/A sky130_fd_sc_hd__clkbuf_2
X_7261_ _7261_/A _7261_/B VGND VGND VPWR VPWR _7263_/A sky130_fd_sc_hd__xnor2_1
X_9000_ _8972_/A _8972_/B _8964_/A VGND VGND VPWR VPWR _9001_/B sky130_fd_sc_hd__o21ba_1
X_6212_ _6294_/A _6212_/B VGND VGND VPWR VPWR _6304_/A sky130_fd_sc_hd__xnor2_2
X_7192_ _7392_/B _7192_/B VGND VGND VPWR VPWR _7195_/A sky130_fd_sc_hd__xnor2_1
X_6143_ _7118_/A _6143_/B VGND VGND VPWR VPWR _6145_/A sky130_fd_sc_hd__and2_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _9171_/Q VGND VGND VPWR VPWR _7327_/A sky130_fd_sc_hd__clkbuf_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _4891_/A _5093_/A _4980_/A VGND VGND VPWR VPWR _5025_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6976_ _7079_/A _6976_/B VGND VGND VPWR VPWR _6978_/C sky130_fd_sc_hd__nor2_1
X_8715_ _8773_/B _8715_/B VGND VGND VPWR VPWR _9102_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5927_ _7096_/A _7627_/A VGND VGND VPWR VPWR _5928_/B sky130_fd_sc_hd__nand2_1
X_8646_ _8568_/A _9025_/B _8569_/A _8567_/B VGND VGND VPWR VPWR _8709_/B sky130_fd_sc_hd__a31oi_2
X_5858_ _5858_/A _5858_/B _5858_/C VGND VGND VPWR VPWR _5858_/X sky130_fd_sc_hd__and3_1
X_5789_ _9193_/Q VGND VGND VPWR VPWR _6235_/A sky130_fd_sc_hd__buf_2
X_8577_ _8504_/B _8513_/Y _8575_/X _8648_/B VGND VGND VPWR VPWR _8579_/A sky130_fd_sc_hd__o211a_1
X_4809_ _4836_/A _4808_/X _5653_/B VGND VGND VPWR VPWR _4810_/A sky130_fd_sc_hd__mux2_1
X_7528_ _7528_/A _7384_/B VGND VGND VPWR VPWR _7528_/X sky130_fd_sc_hd__or2b_1
X_7459_ _8036_/B _8175_/B _7959_/A _7459_/D VGND VGND VPWR VPWR _7460_/B sky130_fd_sc_hd__and4_1
XFILLER_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9129_ _9219_/CLK _9129_/D VGND VGND VPWR VPWR _9129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6830_ _6830_/A _6830_/B VGND VGND VPWR VPWR _6882_/B sky130_fd_sc_hd__xnor2_4
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6761_ _7583_/A _6927_/C _6361_/D _7435_/A VGND VGND VPWR VPWR _6762_/B sky130_fd_sc_hd__a22oi_1
XFILLER_23_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8500_ _8501_/A _8501_/B _8501_/C VGND VGND VPWR VPWR _8500_/Y sky130_fd_sc_hd__o21ai_1
X_5712_ _4636_/A _5711_/X _5712_/S VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__mux2_1
X_6692_ _6691_/A _6691_/B _6691_/C VGND VGND VPWR VPWR _6814_/C sky130_fd_sc_hd__a21oi_4
X_8431_ _8831_/B VGND VGND VPWR VPWR _8891_/B sky130_fd_sc_hd__buf_2
X_5643_ _4573_/X _4637_/A _4643_/A VGND VGND VPWR VPWR _5643_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8362_ _8252_/A _8252_/B _8361_/X VGND VGND VPWR VPWR _8482_/B sky130_fd_sc_hd__a21bo_1
X_5574_ _5433_/A _5573_/X _5671_/S VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
X_7313_ _7203_/A _7313_/B VGND VGND VPWR VPWR _7313_/X sky130_fd_sc_hd__and2b_1
X_8293_ _8530_/A _8466_/A _8542_/A _8542_/B VGND VGND VPWR VPWR _8294_/B sky130_fd_sc_hd__and4_1
XFILLER_104_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7244_ _7244_/A _7244_/B VGND VGND VPWR VPWR _7245_/B sky130_fd_sc_hd__nor2_1
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7175_ _7176_/B _7287_/A _7176_/A VGND VGND VPWR VPWR _7177_/B sky130_fd_sc_hd__o21a_1
XFILLER_105_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6126_ _6126_/A _6126_/B _6049_/C _6125_/A VGND VGND VPWR VPWR _6126_/X sky130_fd_sc_hd__or4bb_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6057_ _6702_/A VGND VGND VPWR VPWR _7037_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5008_ _5007_/A _5044_/A _5006_/X _5007_/Y VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__a31o_1
XFILLER_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _6959_/A _6959_/B VGND VGND VPWR VPWR _7064_/A sky130_fd_sc_hd__nand2_1
X_8629_ _8628_/B _8697_/B _8628_/A VGND VGND VPWR VPWR _8631_/C sky130_fd_sc_hd__a21oi_1
XFILLER_22_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A VGND VGND VPWR VPWR _9221_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5290_ _4847_/X _5430_/A _5288_/X _5289_/X _5151_/A VGND VGND VPWR VPWR _5290_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8980_ _8980_/A _8980_/B VGND VGND VPWR VPWR _8982_/A sky130_fd_sc_hd__xnor2_1
X_7931_ _7932_/A _7932_/B VGND VGND VPWR VPWR _7933_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7862_ _7861_/A _7861_/B _7861_/C VGND VGND VPWR VPWR _7952_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _6940_/A _6940_/B _6940_/C _6940_/D VGND VGND VPWR VPWR _6813_/X sky130_fd_sc_hd__or4_2
X_7793_ _7793_/A _7795_/B _7793_/C VGND VGND VPWR VPWR _7794_/B sky130_fd_sc_hd__nand3_2
X_6744_ _6744_/A _6744_/B VGND VGND VPWR VPWR _6745_/B sky130_fd_sc_hd__xor2_2
X_6675_ _6675_/A _6675_/B _6675_/C VGND VGND VPWR VPWR _6689_/B sky130_fd_sc_hd__nand3_1
X_8414_ _8414_/A _8414_/B VGND VGND VPWR VPWR _8416_/A sky130_fd_sc_hd__nor2_1
X_5626_ _5534_/X _5625_/X _5673_/S VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8345_ _8345_/A VGND VGND VPWR VPWR _8358_/A sky130_fd_sc_hd__inv_2
X_5557_ _5557_/A VGND VGND VPWR VPWR _5754_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8276_ _8792_/D VGND VGND VPWR VPWR _8450_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5488_ _5142_/X _5212_/A _5368_/A VGND VGND VPWR VPWR _5488_/Y sky130_fd_sc_hd__a21oi_1
X_7227_ _7225_/Y _7335_/A _7327_/B _9204_/Q VGND VGND VPWR VPWR _7342_/A sky130_fd_sc_hd__and4bb_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7158_ _7159_/A _7159_/B VGND VGND VPWR VPWR _7160_/A sky130_fd_sc_hd__nor2_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6109_ _7194_/A VGND VGND VPWR VPWR _6875_/A sky130_fd_sc_hd__clkbuf_2
X_7089_ _7088_/A _7088_/B _7088_/C VGND VGND VPWR VPWR _7215_/A sky130_fd_sc_hd__a21oi_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4790_ _5002_/A VGND VGND VPWR VPWR _5214_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 _9135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _5482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6460_ _6512_/A _6512_/B _6546_/A VGND VGND VPWR VPWR _6460_/X sky130_fd_sc_hd__and3_1
X_6391_ _9206_/Q VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5411_ _4667_/A _5630_/A _5408_/X _5409_/Y _5410_/X VGND VGND VPWR VPWR _5411_/X
+ sky130_fd_sc_hd__a221o_1
X_8130_ _8231_/B _8130_/B VGND VGND VPWR VPWR _9095_/D sky130_fd_sc_hd__nor2_1
X_5342_ _4570_/A _5404_/A _5340_/Y _5341_/X _5251_/A VGND VGND VPWR VPWR _5342_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8061_ _8062_/A _8062_/B VGND VGND VPWR VPWR _8063_/A sky130_fd_sc_hd__nand2_1
X_7012_ _7110_/A _7110_/B VGND VGND VPWR VPWR _7013_/C sky130_fd_sc_hd__xnor2_1
X_5273_ _5607_/A VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__buf_2
XFILLER_101_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8963_ _8963_/A _8963_/B _8961_/X VGND VGND VPWR VPWR _8963_/X sky130_fd_sc_hd__or3b_1
X_8894_ _8989_/A _8975_/A VGND VGND VPWR VPWR _8895_/B sky130_fd_sc_hd__nand2_1
X_7914_ _7813_/A _7813_/B _7817_/B VGND VGND VPWR VPWR _7914_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7845_ _7845_/A _7763_/A VGND VGND VPWR VPWR _7861_/B sky130_fd_sc_hd__or2b_1
XFILLER_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7776_ _7656_/B _7776_/B VGND VGND VPWR VPWR _7776_/X sky130_fd_sc_hd__and2b_1
X_4988_ _9126_/Q _9118_/Q VGND VGND VPWR VPWR _4989_/B sky130_fd_sc_hd__or2_1
X_6727_ _7706_/D VGND VGND VPWR VPWR _8720_/A sky130_fd_sc_hd__clkbuf_2
X_6658_ _6658_/A _6599_/A VGND VGND VPWR VPWR _6675_/A sky130_fd_sc_hd__or2b_1
X_5609_ _5149_/X _5122_/A _5607_/Y _5608_/X _5151_/X VGND VGND VPWR VPWR _5609_/X
+ sky130_fd_sc_hd__a221o_1
X_8328_ _8328_/A _8328_/B VGND VGND VPWR VPWR _8336_/B sky130_fd_sc_hd__nand2_1
X_6589_ _6313_/B _7938_/A _7610_/D _6313_/A VGND VGND VPWR VPWR _6591_/A sky130_fd_sc_hd__a22oi_2
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8259_ _8587_/B VGND VGND VPWR VPWR _8832_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput27 A[4] VGND VGND VPWR VPWR _9166_/D sky130_fd_sc_hd__clkbuf_1
Xinput16 A[23] VGND VGND VPWR VPWR _9185_/D sky130_fd_sc_hd__clkbuf_1
Xinput49 B[24] VGND VGND VPWR VPWR _9217_/D sky130_fd_sc_hd__clkbuf_1
Xinput38 B[14] VGND VGND VPWR VPWR _9207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5960_ _7627_/A VGND VGND VPWR VPWR _8071_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4911_ _4950_/B VGND VGND VPWR VPWR _4957_/B sky130_fd_sc_hd__clkbuf_2
X_5891_ _7645_/A _6359_/A _6828_/A _7647_/A VGND VGND VPWR VPWR _5892_/B sky130_fd_sc_hd__a22oi_2
X_7630_ _7490_/B _7754_/A _7629_/Y VGND VGND VPWR VPWR _7633_/A sky130_fd_sc_hd__a21oi_1
XFILLER_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4842_ _4842_/A _4842_/B VGND VGND VPWR VPWR _4845_/A sky130_fd_sc_hd__or2_1
X_7561_ _7561_/A _7561_/B VGND VGND VPWR VPWR _7563_/A sky130_fd_sc_hd__nor2_1
X_4773_ _4929_/A _4924_/A VGND VGND VPWR VPWR _4773_/Y sky130_fd_sc_hd__nor2_1
X_7492_ _7492_/A _7492_/B VGND VGND VPWR VPWR _7493_/B sky130_fd_sc_hd__xnor2_1
X_6512_ _6512_/A _6512_/B _6546_/A VGND VGND VPWR VPWR _6546_/B sky130_fd_sc_hd__nand3_1
X_6443_ _7016_/A _6590_/B _7706_/A _7465_/A VGND VGND VPWR VPWR _6444_/B sky130_fd_sc_hd__and4_1
X_6374_ _6375_/A _6466_/A _6375_/C VGND VGND VPWR VPWR _6376_/A sky130_fd_sc_hd__a21oi_1
X_9162_ _9220_/CLK input1/X VGND VGND VPWR VPWR _9162_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8113_ _8005_/A _8005_/B _8008_/B VGND VGND VPWR VPWR _8114_/B sky130_fd_sc_hd__o21ba_1
X_5325_ _5213_/X _5212_/X _4723_/X VGND VGND VPWR VPWR _5325_/Y sky130_fd_sc_hd__a21oi_1
X_9093_ _9212_/CLK _9093_/D VGND VGND VPWR VPWR _9093_/Q sky130_fd_sc_hd__dfxtp_1
X_8044_ _8220_/A _8044_/B VGND VGND VPWR VPWR _8045_/B sky130_fd_sc_hd__nand2_1
X_5256_ _5618_/A _5430_/A _5254_/X _5255_/X _4566_/A VGND VGND VPWR VPWR _5256_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _5187_/A VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__clkbuf_2
X_8946_ _8947_/A _8947_/B VGND VGND VPWR VPWR _8948_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8877_ _8878_/A _8878_/B _8878_/C VGND VGND VPWR VPWR _8921_/A sky130_fd_sc_hd__o21ai_1
XFILLER_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7828_ _7828_/A _7828_/B _7828_/C VGND VGND VPWR VPWR _7829_/B sky130_fd_sc_hd__nor3_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7759_ _7759_/A _7759_/B VGND VGND VPWR VPWR _7761_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6090_/A _6090_/B _6090_/C VGND VGND VPWR VPWR _6104_/C sky130_fd_sc_hd__nand3_2
X_5110_ _5676_/B _5108_/X _5109_/X _5506_/A VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__o211a_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A VGND VGND VPWR VPWR _5043_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8800_ _8800_/A _8800_/B VGND VGND VPWR VPWR _8865_/B sky130_fd_sc_hd__nand2_1
X_8731_ _8805_/A _8731_/B VGND VGND VPWR VPWR _8744_/A sky130_fd_sc_hd__xor2_1
XFILLER_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6992_ _7075_/A _7174_/B VGND VGND VPWR VPWR _7058_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5943_ _7299_/A VGND VGND VPWR VPWR _7531_/A sky130_fd_sc_hd__clkbuf_2
X_8662_ _8662_/A _8662_/B VGND VGND VPWR VPWR _8671_/A sky130_fd_sc_hd__or2_1
X_5874_ _6825_/B VGND VGND VPWR VPWR _6858_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8593_ _8688_/A _8593_/B VGND VGND VPWR VPWR _8628_/A sky130_fd_sc_hd__nor2_1
X_7613_ _7470_/A _7469_/A _7469_/B VGND VGND VPWR VPWR _7614_/B sky130_fd_sc_hd__o21ba_1
XFILLER_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4825_ _4928_/A VGND VGND VPWR VPWR _4845_/B sky130_fd_sc_hd__clkbuf_2
X_7544_ _7544_/A _7544_/B _7544_/C VGND VGND VPWR VPWR _7553_/A sky130_fd_sc_hd__and3_1
X_4756_ _4824_/A VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7475_ _7474_/A _7474_/B _7474_/C VGND VGND VPWR VPWR _7475_/X sky130_fd_sc_hd__a21o_4
X_4687_ _9111_/Q VGND VGND VPWR VPWR _4687_/X sky130_fd_sc_hd__clkbuf_2
X_6426_ _7083_/B VGND VGND VPWR VPWR _7419_/B sky130_fd_sc_hd__clkbuf_2
X_9214_ _9214_/CLK _9214_/D VGND VGND VPWR VPWR _9214_/Q sky130_fd_sc_hd__dfxtp_2
X_6357_ _8086_/A VGND VGND VPWR VPWR _8517_/A sky130_fd_sc_hd__clkbuf_4
X_9145_ _9214_/CLK _9145_/D VGND VGND VPWR VPWR _9145_/Q sky130_fd_sc_hd__dfxtp_1
X_5308_ _5697_/S VGND VGND VPWR VPWR _5428_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9076_ _9214_/CLK _9076_/D VGND VGND VPWR VPWR _9076_/Q sky130_fd_sc_hd__dfxtp_1
X_6288_ _6288_/A _6288_/B _6288_/C VGND VGND VPWR VPWR _6288_/X sky130_fd_sc_hd__and3_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8027_ _7918_/A _8949_/B _7919_/A _7917_/B VGND VGND VPWR VPWR _8132_/A sky130_fd_sc_hd__a31o_1
X_5239_ _5206_/X _5237_/X _5281_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8929_ _8929_/A _8929_/B _8929_/C VGND VGND VPWR VPWR _8979_/B sky130_fd_sc_hd__and3_1
XFILLER_44_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4610_ _5735_/S VGND VGND VPWR VPWR _5691_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5590_ _5258_/A _5116_/A _5588_/X _5589_/Y _4598_/A VGND VGND VPWR VPWR _5590_/X
+ sky130_fd_sc_hd__a221o_1
X_4541_ _4541_/A VGND VGND VPWR VPWR _4541_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7260_ _7260_/A _7260_/B VGND VGND VPWR VPWR _7261_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6211_ _6211_/A _6211_/B VGND VGND VPWR VPWR _6212_/B sky130_fd_sc_hd__or2_1
X_7191_ _7094_/A _7097_/B _7094_/B VGND VGND VPWR VPWR _7192_/B sky130_fd_sc_hd__o21ba_1
X_6142_ _9171_/Q VGND VGND VPWR VPWR _6143_/B sky130_fd_sc_hd__buf_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6073_ _6530_/B VGND VGND VPWR VPWR _6313_/B sky130_fd_sc_hd__clkbuf_2
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _4538_/A _4940_/C _5022_/X _5023_/X _4739_/X VGND VGND VPWR VPWR _5024_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6975_ _6405_/B _6825_/C _7822_/D _7293_/A VGND VGND VPWR VPWR _6976_/B sky130_fd_sc_hd__a22oi_1
X_5926_ _7869_/A VGND VGND VPWR VPWR _7627_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8714_ _8770_/A _8714_/B VGND VGND VPWR VPWR _8715_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8645_ _8645_/A _8645_/B VGND VGND VPWR VPWR _8709_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5857_ _6974_/A _7365_/A _5810_/X _5809_/X _5940_/A VGND VGND VPWR VPWR _5858_/C
+ sky130_fd_sc_hd__a32o_1
X_8576_ _8496_/B _8499_/B _8573_/X _8648_/A VGND VGND VPWR VPWR _8648_/B sky130_fd_sc_hd__o211ai_2
X_4808_ _5510_/A _4760_/X _4807_/X VGND VGND VPWR VPWR _4808_/X sky130_fd_sc_hd__o21a_1
X_5788_ _6974_/B VGND VGND VPWR VPWR _7201_/A sky130_fd_sc_hd__buf_2
X_7527_ _7527_/A _7559_/B _7527_/C _7665_/A VGND VGND VPWR VPWR _7665_/B sky130_fd_sc_hd__nor4_2
X_4739_ _4739_/A VGND VGND VPWR VPWR _4739_/X sky130_fd_sc_hd__clkbuf_2
X_7458_ _8175_/B _7959_/A _8084_/A _8036_/B VGND VGND VPWR VPWR _7460_/A sky130_fd_sc_hd__a22oi_1
XFILLER_79_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6409_ _6409_/A _6485_/A VGND VGND VPWR VPWR _6410_/B sky130_fd_sc_hd__xnor2_1
X_7389_ _7389_/A _9215_/Q VGND VGND VPWR VPWR _7397_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9128_ _9223_/CLK hold13/X VGND VGND VPWR VPWR _9128_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9059_ _9059_/A _9059_/B _9062_/A VGND VGND VPWR VPWR _9059_/X sky130_fd_sc_hd__or3_1
XFILLER_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6760_ _6760_/A VGND VGND VPWR VPWR _7583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5711_ _5460_/A _5170_/X _5709_/X _5710_/Y VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__a22o_1
X_6691_ _6691_/A _6691_/B _6691_/C VGND VGND VPWR VPWR _6814_/B sky130_fd_sc_hd__and3_1
X_8430_ _8430_/A _8430_/B VGND VGND VPWR VPWR _9098_/D sky130_fd_sc_hd__xnor2_1
X_5642_ _5314_/A _4874_/S _5640_/X _5641_/Y _5382_/X VGND VGND VPWR VPWR _5642_/X
+ sky130_fd_sc_hd__a221o_1
X_8361_ _8361_/A _8251_/A VGND VGND VPWR VPWR _8361_/X sky130_fd_sc_hd__or2b_1
X_5573_ _4635_/A _5572_/X _5670_/S VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__mux2_1
X_7312_ _7312_/A _7312_/B VGND VGND VPWR VPWR _7316_/A sky130_fd_sc_hd__xnor2_1
X_8292_ _8607_/B VGND VGND VPWR VPWR _8542_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7243_ _7349_/A _9200_/Q _9176_/Q _9177_/Q VGND VGND VPWR VPWR _7244_/B sky130_fd_sc_hd__and4_1
X_7174_ _7174_/A _7174_/B VGND VGND VPWR VPWR _7176_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6125_ _6125_/A _6125_/B VGND VGND VPWR VPWR _6128_/A sky130_fd_sc_hd__xnor2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6056_ _7006_/B VGND VGND VPWR VPWR _6223_/B sky130_fd_sc_hd__buf_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5007_ _5007_/A _5007_/B VGND VGND VPWR VPWR _5007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6958_ _6956_/Y _6955_/B _6957_/X VGND VGND VPWR VPWR _7065_/A sky130_fd_sc_hd__a21bo_1
X_6889_ _9198_/Q _7241_/B VGND VGND VPWR VPWR _6891_/A sky130_fd_sc_hd__and2_1
X_5909_ _9168_/Q VGND VGND VPWR VPWR _6232_/A sky130_fd_sc_hd__buf_2
X_8628_ _8628_/A _8628_/B _8697_/B VGND VGND VPWR VPWR _8694_/A sky130_fd_sc_hd__and3_1
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8559_ _8559_/A _8559_/B _8635_/B VGND VGND VPWR VPWR _8631_/A sky130_fd_sc_hd__or3_2
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7930_ _8032_/A _8044_/B VGND VGND VPWR VPWR _7932_/B sky130_fd_sc_hd__and2_1
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7861_ _7861_/A _7861_/B _7861_/C VGND VGND VPWR VPWR _7863_/A sky130_fd_sc_hd__nand3_1
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6812_ _6940_/A _6940_/B _6940_/C _6940_/D VGND VGND VPWR VPWR _6812_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_90_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7792_ _7793_/A _7795_/B _7793_/C VGND VGND VPWR VPWR _7792_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6743_ _6743_/A _6845_/C VGND VGND VPWR VPWR _6744_/B sky130_fd_sc_hd__xnor2_2
X_6674_ _6774_/A _6774_/B VGND VGND VPWR VPWR _6675_/C sky130_fd_sc_hd__xnor2_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8413_ _8412_/A _8412_/B _8411_/Y VGND VGND VPWR VPWR _8414_/B sky130_fd_sc_hd__o21ba_1
X_5625_ _5509_/A _4769_/A _5623_/X _5624_/Y VGND VGND VPWR VPWR _5625_/X sky130_fd_sc_hd__a22o_1
X_8344_ _8344_/A _8470_/B VGND VGND VPWR VPWR _8345_/A sky130_fd_sc_hd__nor2_1
X_5556_ _5534_/X _5510_/X _5511_/X _5554_/X _5555_/X VGND VGND VPWR VPWR _9141_/D
+ sky130_fd_sc_hd__o221a_4
X_8275_ _8452_/A _8978_/A _8974_/A _8371_/A VGND VGND VPWR VPWR _8278_/A sky130_fd_sc_hd__a22oi_1
X_5487_ _5149_/X _9081_/Q _5485_/Y _5486_/X _5151_/X VGND VGND VPWR VPWR _5487_/X
+ sky130_fd_sc_hd__a221o_1
X_7226_ _9202_/Q _9203_/Q _9173_/Q _9174_/Q VGND VGND VPWR VPWR _7335_/A sky130_fd_sc_hd__and4_1
X_7157_ _7237_/B _7157_/B VGND VGND VPWR VPWR _7159_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A _6108_/B VGND VGND VPWR VPWR _6108_/X sky130_fd_sc_hd__and2_1
X_7088_ _7088_/A _7088_/B _7088_/C VGND VGND VPWR VPWR _7102_/B sky130_fd_sc_hd__and3_1
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6039_ _6037_/A _6037_/Y _6035_/X _6036_/Y VGND VGND VPWR VPWR _6041_/C sky130_fd_sc_hd__a211o_1
XFILLER_100_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_19 _9135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6390_ _7604_/C VGND VGND VPWR VPWR _7959_/A sky130_fd_sc_hd__buf_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5410_ _5410_/A VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5341_ _4849_/A _5370_/A _5146_/X _5316_/A _4783_/X VGND VGND VPWR VPWR _5341_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8060_ _8060_/A _8060_/B VGND VGND VPWR VPWR _8062_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7011_ _7011_/A _7109_/A VGND VGND VPWR VPWR _7110_/B sky130_fd_sc_hd__xnor2_1
X_5272_ _9084_/Q VGND VGND VPWR VPWR _5607_/A sky130_fd_sc_hd__inv_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8962_ _8963_/A _8963_/B _8961_/X VGND VGND VPWR VPWR _8964_/A sky130_fd_sc_hd__o21ba_1
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7913_ _7804_/A _8949_/B _7805_/A _7803_/B VGND VGND VPWR VPWR _8016_/A sky130_fd_sc_hd__a31o_1
XFILLER_102_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8893_ _8842_/X _8925_/A _8892_/Y VGND VGND VPWR VPWR _8895_/A sky130_fd_sc_hd__a21oi_1
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7844_ _7739_/A _7739_/B _7843_/X VGND VGND VPWR VPWR _7920_/A sky130_fd_sc_hd__a21oi_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7775_ _7865_/A _7865_/B VGND VGND VPWR VPWR _7895_/A sky130_fd_sc_hd__xnor2_4
X_6726_ _9209_/Q VGND VGND VPWR VPWR _7706_/D sky130_fd_sc_hd__clkbuf_2
X_4987_ _9126_/Q _9118_/Q VGND VGND VPWR VPWR _5032_/A sky130_fd_sc_hd__nand2_1
X_6657_ _6646_/A _6646_/B _6656_/Y VGND VGND VPWR VPWR _6750_/A sky130_fd_sc_hd__o21a_1
X_6588_ _7116_/D VGND VGND VPWR VPWR _7610_/D sky130_fd_sc_hd__buf_2
X_5608_ _5371_/A _5208_/A _4660_/A _5210_/A _4571_/A VGND VGND VPWR VPWR _5608_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A VGND VGND VPWR VPWR _9223_/CLK sky130_fd_sc_hd__clkbuf_2
X_8327_ _8223_/C _8224_/B _8324_/Y _8325_/X VGND VGND VPWR VPWR _8328_/B sky130_fd_sc_hd__o211ai_2
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5539_ _4634_/A _5208_/A _5538_/X _4593_/A VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__a211o_1
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8258_ _8258_/A VGND VGND VPWR VPWR _8365_/A sky130_fd_sc_hd__inv_2
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8189_ _8290_/A _8190_/C _8607_/B _8190_/A VGND VGND VPWR VPWR _8191_/A sky130_fd_sc_hd__a22oi_1
X_7209_ _7209_/A _7209_/B VGND VGND VPWR VPWR _7321_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 A[24] VGND VGND VPWR VPWR _9186_/D sky130_fd_sc_hd__clkbuf_1
Xinput28 A[5] VGND VGND VPWR VPWR _9167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 B[15] VGND VGND VPWR VPWR _9208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5890_ _5922_/A VGND VGND VPWR VPWR _6828_/A sky130_fd_sc_hd__clkbuf_2
X_4910_ _5044_/A VGND VGND VPWR VPWR _4950_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4841_ _4841_/A VGND VGND VPWR VPWR _5249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7560_ _7559_/A _7559_/B _7558_/Y VGND VGND VPWR VPWR _7561_/B sky130_fd_sc_hd__o21ba_1
XFILLER_33_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4772_ _5181_/A VGND VGND VPWR VPWR _5403_/A sky130_fd_sc_hd__clkbuf_2
X_7491_ _7487_/Y _7629_/A _7490_/Y VGND VGND VPWR VPWR _7492_/B sky130_fd_sc_hd__a21oi_2
X_6511_ _6622_/A _6622_/B VGND VGND VPWR VPWR _6548_/A sky130_fd_sc_hd__xnor2_1
X_6442_ _7131_/C VGND VGND VPWR VPWR _7465_/A sky130_fd_sc_hd__clkbuf_2
X_9161_ _9224_/CLK _9161_/D VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
X_8112_ _8112_/A _8211_/B VGND VGND VPWR VPWR _8114_/A sky130_fd_sc_hd__nand2_1
X_6373_ _6288_/A _6288_/B _6288_/C VGND VGND VPWR VPWR _6375_/C sky130_fd_sc_hd__a21bo_1
X_5324_ _5164_/A _5604_/A _5322_/X _5323_/Y _4923_/A VGND VGND VPWR VPWR _5324_/X
+ sky130_fd_sc_hd__a221o_1
X_9092_ _9212_/CLK _9092_/D VGND VGND VPWR VPWR _9092_/Q sky130_fd_sc_hd__dfxtp_1
X_8043_ _8215_/B _8043_/B VGND VGND VPWR VPWR _8045_/A sky130_fd_sc_hd__xnor2_1
X_5255_ _5149_/A _9073_/Q _5151_/A VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__a21o_1
X_5186_ _5020_/X _5124_/X _5182_/X _5185_/Y _4697_/A VGND VGND VPWR VPWR _5186_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8945_ _8945_/A _8945_/B VGND VGND VPWR VPWR _8947_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8876_ _8876_/A _8876_/B VGND VGND VPWR VPWR _8878_/C sky130_fd_sc_hd__xor2_1
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7827_ _7828_/A _7828_/B _7828_/C VGND VGND VPWR VPWR _7946_/B sky130_fd_sc_hd__o21a_1
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7758_ _7873_/A _8150_/D VGND VGND VPWR VPWR _7759_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7689_ _7689_/A _7804_/B VGND VGND VPWR VPWR _7690_/B sky130_fd_sc_hd__nand2_1
X_6709_ _6709_/A _6709_/B VGND VGND VPWR VPWR _6710_/C sky130_fd_sc_hd__xnor2_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6991_ _6869_/B _6878_/B _6988_/X _7174_/A VGND VGND VPWR VPWR _7174_/B sky130_fd_sc_hd__a211oi_1
X_8730_ _8671_/A _8671_/B _8670_/B VGND VGND VPWR VPWR _8731_/B sky130_fd_sc_hd__a21o_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5942_ _7189_/C VGND VGND VPWR VPWR _7299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8661_ _8661_/A _8661_/B _8662_/B VGND VGND VPWR VPWR _8672_/A sky130_fd_sc_hd__or3_1
X_5873_ _5985_/A VGND VGND VPWR VPWR _6825_/B sky130_fd_sc_hd__buf_2
X_8592_ _8591_/B _8592_/B VGND VGND VPWR VPWR _8593_/B sky130_fd_sc_hd__and2b_1
X_7612_ _7612_/A _7612_/B VGND VGND VPWR VPWR _7742_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4824_ _4824_/A _4828_/C VGND VGND VPWR VPWR _4943_/A sky130_fd_sc_hd__nand2_4
X_4755_ _4828_/B VGND VGND VPWR VPWR _4824_/A sky130_fd_sc_hd__buf_2
X_7543_ _7543_/A _7543_/B VGND VGND VPWR VPWR _7544_/C sky130_fd_sc_hd__xnor2_1
X_9213_ _9213_/CLK _9213_/D VGND VGND VPWR VPWR _9213_/Q sky130_fd_sc_hd__dfxtp_2
X_7474_ _7474_/A _7474_/B _7474_/C VGND VGND VPWR VPWR _7474_/Y sky130_fd_sc_hd__nand3_2
X_4686_ _4982_/A VGND VGND VPWR VPWR _5510_/A sky130_fd_sc_hd__clkbuf_2
X_6425_ _6425_/A _6425_/B VGND VGND VPWR VPWR _6430_/A sky130_fd_sc_hd__nor2_1
X_6356_ _7847_/A VGND VGND VPWR VPWR _8086_/A sky130_fd_sc_hd__clkbuf_2
X_9144_ _9199_/CLK _9144_/D VGND VGND VPWR VPWR _9144_/Q sky130_fd_sc_hd__dfxtp_1
X_9075_ _9214_/CLK _9075_/D VGND VGND VPWR VPWR _9075_/Q sky130_fd_sc_hd__dfxtp_4
X_5307_ _5117_/X _5305_/X _5427_/S VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8026_ _8128_/B VGND VGND VPWR VPWR _8026_/Y sky130_fd_sc_hd__inv_2
X_6287_ _6288_/B _6288_/C _6288_/A VGND VGND VPWR VPWR _6287_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5238_ _5740_/S VGND VGND VPWR VPWR _5281_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5169_ _5169_/A VGND VGND VPWR VPWR _5414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8928_ _8929_/A _8929_/B _8929_/C VGND VGND VPWR VPWR _8930_/A sky130_fd_sc_hd__a21oi_1
XFILLER_83_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8859_ _8859_/A _8859_/B VGND VGND VPWR VPWR _8860_/B sky130_fd_sc_hd__or2_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4540_ _5391_/A VGND VGND VPWR VPWR _4541_/A sky130_fd_sc_hd__clkbuf_2
X_6210_ _6210_/A _6210_/B _6210_/C VGND VGND VPWR VPWR _6211_/B sky130_fd_sc_hd__and3_1
X_7190_ _7190_/A _7190_/B VGND VGND VPWR VPWR _7392_/B sky130_fd_sc_hd__nor2_1
X_6141_ _7365_/A VGND VGND VPWR VPWR _7118_/A sky130_fd_sc_hd__clkbuf_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _7083_/B VGND VGND VPWR VPWR _6754_/B sky130_fd_sc_hd__clkbuf_2
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5305_/S _4932_/X _5696_/S VGND VGND VPWR VPWR _5023_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6974_ _6974_/A _6974_/B _9208_/Q _7307_/D VGND VGND VPWR VPWR _7079_/A sky130_fd_sc_hd__and4_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5925_ _7131_/A VGND VGND VPWR VPWR _7869_/A sky130_fd_sc_hd__clkbuf_4
X_8713_ _8648_/A _8648_/B _8649_/A VGND VGND VPWR VPWR _8770_/A sky130_fd_sc_hd__a21o_1
XFILLER_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8644_ _8644_/A _8644_/B VGND VGND VPWR VPWR _8645_/B sky130_fd_sc_hd__or2_1
X_5856_ _6014_/A VGND VGND VPWR VPWR _6974_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ _4535_/A _4764_/X _4804_/X _4806_/Y _9112_/Q VGND VGND VPWR VPWR _4807_/X
+ sky130_fd_sc_hd__a221o_1
X_8575_ _8573_/X _8648_/A _8496_/B _8499_/B VGND VGND VPWR VPWR _8575_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5787_ _9166_/Q VGND VGND VPWR VPWR _6974_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7526_ _7527_/A _7559_/B _7527_/C _7665_/A VGND VGND VPWR VPWR _7526_/X sky130_fd_sc_hd__o22a_1
X_4738_ _4889_/A _4698_/X _4736_/Y _4737_/X VGND VGND VPWR VPWR _4738_/X sky130_fd_sc_hd__a211o_1
X_7457_ _7457_/A VGND VGND VPWR VPWR _8036_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4669_ _9090_/Q VGND VGND VPWR VPWR _5393_/A sky130_fd_sc_hd__buf_2
X_6408_ _6363_/A _6362_/A _6362_/B VGND VGND VPWR VPWR _6485_/A sky130_fd_sc_hd__o21ba_1
X_9127_ _9222_/CLK hold6/X VGND VGND VPWR VPWR _9127_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7388_ _7277_/D _7277_/Y _7385_/Y _7386_/X VGND VGND VPWR VPWR _7539_/C sky130_fd_sc_hd__o211ai_4
X_6339_ _7083_/B _7307_/A _6680_/A _6680_/B VGND VGND VPWR VPWR _6340_/B sky130_fd_sc_hd__and4_1
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9058_ _9058_/A VGND VGND VPWR VPWR _9071_/D sky130_fd_sc_hd__clkbuf_1
X_8009_ _7897_/A _8009_/B VGND VGND VPWR VPWR _8009_/X sky130_fd_sc_hd__and2b_2
XFILLER_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5710_ _5621_/X _5132_/X _4642_/A VGND VGND VPWR VPWR _5710_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6690_ _6690_/A _6810_/B VGND VGND VPWR VPWR _6691_/C sky130_fd_sc_hd__nand2_1
X_5641_ _5450_/A _4600_/A _5367_/X VGND VGND VPWR VPWR _5641_/Y sky130_fd_sc_hd__a21oi_1
X_8360_ _8481_/A _8481_/B VGND VGND VPWR VPWR _8363_/A sky130_fd_sc_hd__xnor2_1
X_5572_ _4587_/X _5571_/Y _5572_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
X_8291_ _8595_/A _8664_/A _8664_/B _8530_/A VGND VGND VPWR VPWR _8294_/A sky130_fd_sc_hd__a22oi_1
X_7311_ _7311_/A _7441_/B VGND VGND VPWR VPWR _7312_/B sky130_fd_sc_hd__xnor2_1
X_7242_ _7019_/B _7131_/D _9177_/Q _7348_/A VGND VGND VPWR VPWR _7244_/A sky130_fd_sc_hd__a22oi_1
X_7173_ _7172_/A _7172_/B _7172_/C VGND VGND VPWR VPWR _7287_/A sky130_fd_sc_hd__a21oi_2
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6124_ _6221_/B _6124_/B VGND VGND VPWR VPWR _6125_/B sky130_fd_sc_hd__xnor2_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A VGND VGND VPWR VPWR _7006_/B sky130_fd_sc_hd__clkbuf_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4943_/A _5004_/Y _5005_/X _4706_/S VGND VGND VPWR VPWR _5006_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6957_ _6957_/A _6957_/B VGND VGND VPWR VPWR _6957_/X sky130_fd_sc_hd__or2_1
XFILLER_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6888_ _6998_/B _7346_/B _7119_/D _6998_/A VGND VGND VPWR VPWR _6891_/C sky130_fd_sc_hd__a22o_1
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5908_ _6702_/A _5908_/B VGND VGND VPWR VPWR _5987_/B sky130_fd_sc_hd__nand2_1
X_8627_ _8627_/A VGND VGND VPWR VPWR _8697_/B sky130_fd_sc_hd__inv_2
X_5839_ _9197_/Q VGND VGND VPWR VPWR _7253_/B sky130_fd_sc_hd__buf_2
X_8558_ _8478_/B _8480_/X _8555_/Y _8635_/A VGND VGND VPWR VPWR _8635_/B sky130_fd_sc_hd__a211oi_4
X_7509_ _7509_/A _7769_/A VGND VGND VPWR VPWR _7510_/B sky130_fd_sc_hd__nand2_1
X_8489_ _8562_/A _8489_/B VGND VGND VPWR VPWR _8490_/C sky130_fd_sc_hd__nor2_1
XFILLER_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7860_ _7860_/A _7860_/B VGND VGND VPWR VPWR _7861_/C sky130_fd_sc_hd__or2_1
X_6811_ _6810_/A _6810_/B _6810_/C VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__a21oi_4
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7791_ _7791_/A _7791_/B VGND VGND VPWR VPWR _7793_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6742_ _6640_/A _6640_/B _6640_/C VGND VGND VPWR VPWR _6845_/C sky130_fd_sc_hd__a21bo_1
X_6673_ _6673_/A _6773_/A VGND VGND VPWR VPWR _6774_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8412_ _8412_/A _8412_/B _8411_/Y VGND VGND VPWR VPWR _8414_/A sky130_fd_sc_hd__nor3b_1
X_5624_ _4872_/S _5020_/X _4697_/A VGND VGND VPWR VPWR _5624_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8343_ _8343_/A _8470_/A _8343_/C VGND VGND VPWR VPWR _8470_/B sky130_fd_sc_hd__nor3_1
X_5555_ _5555_/A _5604_/B VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__or2_1
XFILLER_104_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8274_ _8844_/C VGND VGND VPWR VPWR _8974_/A sky130_fd_sc_hd__clkbuf_2
X_5486_ _5371_/A _5131_/A _4660_/A _5248_/A _4572_/A VGND VGND VPWR VPWR _5486_/X
+ sky130_fd_sc_hd__o221a_1
X_7225_ _7152_/C _9173_/Q _7019_/C _7152_/A VGND VGND VPWR VPWR _7225_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_104_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7156_ _7044_/A _7043_/A _7043_/B VGND VGND VPWR VPWR _7157_/B sky130_fd_sc_hd__o21ba_1
XFILLER_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6107_/A _6107_/B VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__and2_1
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7087_ _7087_/A _7087_/B VGND VGND VPWR VPWR _7088_/C sky130_fd_sc_hd__xnor2_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6038_ _6035_/X _6036_/Y _6037_/A _6037_/Y VGND VGND VPWR VPWR _6041_/B sky130_fd_sc_hd__o211ai_2
XFILLER_27_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7989_ _7990_/A _7990_/B _7990_/C VGND VGND VPWR VPWR _7991_/A sky130_fd_sc_hd__a21oi_1
XFILLER_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ _9074_/Q _5559_/B VGND VGND VPWR VPWR _5340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5271_ _5271_/A VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7010_ _6897_/A _6896_/B _6896_/A VGND VGND VPWR VPWR _7109_/A sky130_fd_sc_hd__o21ba_1
XFILLER_101_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8961_ _8961_/A _8973_/B VGND VGND VPWR VPWR _8961_/X sky130_fd_sc_hd__xor2_1
XFILLER_95_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7912_ _8639_/B VGND VGND VPWR VPWR _8949_/B sky130_fd_sc_hd__buf_2
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8892_ _8974_/A _9004_/A _8891_/B _8978_/A VGND VGND VPWR VPWR _8892_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7843_ _7738_/B _7843_/B VGND VGND VPWR VPWR _7843_/X sky130_fd_sc_hd__and2b_1
XFILLER_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7774_ _7774_/A _7891_/A VGND VGND VPWR VPWR _7865_/B sky130_fd_sc_hd__and2_2
X_4986_ _4905_/A _4991_/A _4904_/B _4913_/A _4913_/B VGND VGND VPWR VPWR _4994_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6725_ _8190_/C VGND VGND VPWR VPWR _8721_/A sky130_fd_sc_hd__clkbuf_4
X_6656_ _6656_/A _6656_/B VGND VGND VPWR VPWR _6656_/Y sky130_fd_sc_hd__nand2_1
X_6587_ _9177_/Q VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5607_ _5607_/A _5634_/B VGND VGND VPWR VPWR _5607_/Y sky130_fd_sc_hd__nand2_1
X_8326_ _8324_/Y _8325_/X _8223_/C _8224_/B VGND VGND VPWR VPWR _8328_/A sky130_fd_sc_hd__a211o_1
X_5538_ _5618_/A _5124_/A _5536_/Y _5537_/X _4566_/A VGND VGND VPWR VPWR _5538_/X
+ sky130_fd_sc_hd__o221a_1
X_8257_ _8138_/B _8257_/B _8257_/C VGND VGND VPWR VPWR _8258_/A sky130_fd_sc_hd__and3b_1
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5469_ _5214_/X _5634_/A _5467_/X _5468_/Y _5001_/A VGND VGND VPWR VPWR _5469_/X
+ sky130_fd_sc_hd__a221o_1
X_7208_ _7208_/A _7208_/B VGND VGND VPWR VPWR _7209_/B sky130_fd_sc_hd__or2_1
X_8188_ _8087_/A _8089_/B _8087_/B VGND VGND VPWR VPWR _8195_/A sky130_fd_sc_hd__o21ba_1
XFILLER_59_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7139_ _7139_/A _7139_/B _7139_/C VGND VGND VPWR VPWR _7140_/B sky130_fd_sc_hd__nand3_2
XFILLER_59_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 A[25] VGND VGND VPWR VPWR _9187_/D sky130_fd_sc_hd__clkbuf_1
Xinput29 A[6] VGND VGND VPWR VPWR _9168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4840_ _5215_/A VGND VGND VPWR VPWR _4841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6510_ _6508_/X _6637_/A VGND VGND VPWR VPWR _6622_/B sky130_fd_sc_hd__and2b_1
X_4771_ _9106_/Q VGND VGND VPWR VPWR _5181_/A sky130_fd_sc_hd__clkbuf_2
X_7490_ _7490_/A _7490_/B VGND VGND VPWR VPWR _7490_/Y sky130_fd_sc_hd__nor2_1
X_6441_ _9175_/Q VGND VGND VPWR VPWR _7131_/C sky130_fd_sc_hd__clkbuf_2
X_9160_ _9216_/CLK hold15/X VGND VGND VPWR VPWR _9160_/Q sky130_fd_sc_hd__dfxtp_1
X_6372_ _6372_/A _6372_/B _6372_/C VGND VGND VPWR VPWR _6466_/A sky130_fd_sc_hd__or3_1
X_8111_ _8111_/A _8217_/B _8111_/C VGND VGND VPWR VPWR _8211_/B sky130_fd_sc_hd__or3_1
X_5323_ _4598_/A _5246_/Y _4556_/A VGND VGND VPWR VPWR _5323_/Y sky130_fd_sc_hd__a21oi_1
X_9091_ _9212_/CLK _9091_/D VGND VGND VPWR VPWR _9091_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8042_ _7924_/A _7927_/B _7924_/B VGND VGND VPWR VPWR _8043_/B sky130_fd_sc_hd__o21ba_1
X_5254_ _9071_/Q _4580_/X _4676_/C _9070_/Q _5253_/X VGND VGND VPWR VPWR _5254_/X
+ sky130_fd_sc_hd__o221a_1
X_5185_ _4883_/X _5184_/X _4770_/X VGND VGND VPWR VPWR _5185_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8944_ _8944_/A _8897_/A VGND VGND VPWR VPWR _8945_/A sky130_fd_sc_hd__or2b_1
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8875_ _8816_/A _9004_/B _8815_/B _8813_/X VGND VGND VPWR VPWR _8876_/B sky130_fd_sc_hd__a31o_1
X_7826_ _7826_/A _7934_/B VGND VGND VPWR VPWR _7828_/C sky130_fd_sc_hd__xnor2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7757_ _8148_/A VGND VGND VPWR VPWR _8150_/D sky130_fd_sc_hd__buf_2
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4969_ _4922_/X _4968_/Y _4629_/A VGND VGND VPWR VPWR _4969_/X sky130_fd_sc_hd__a21o_1
X_7688_ _7688_/A _7688_/B VGND VGND VPWR VPWR _7690_/A sky130_fd_sc_hd__nor2_1
X_6708_ _6769_/B _6708_/B VGND VGND VPWR VPWR _6709_/B sky130_fd_sc_hd__xnor2_1
X_6639_ _6640_/B _6640_/C _6640_/A VGND VGND VPWR VPWR _6641_/A sky130_fd_sc_hd__a21oi_1
X_8309_ _8165_/B _8168_/C _8306_/X _8307_/Y VGND VGND VPWR VPWR _8412_/A sky130_fd_sc_hd__a211oi_4
XFILLER_3_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6990_ _6988_/X _7174_/A _6869_/B _6878_/B VGND VGND VPWR VPWR _7075_/A sky130_fd_sc_hd__o211a_1
Xclkbuf_4_1_0_clk clkbuf_4_1_0_clk/A VGND VGND VPWR VPWR _9218_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5941_ _7093_/B VGND VGND VPWR VPWR _7189_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5872_ _7506_/B VGND VGND VPWR VPWR _7647_/A sky130_fd_sc_hd__buf_4
X_8660_ _8716_/A _8832_/B _8660_/C VGND VGND VPWR VPWR _8726_/A sky130_fd_sc_hd__and3_1
X_8591_ _8592_/B _8591_/B VGND VGND VPWR VPWR _8688_/A sky130_fd_sc_hd__and2b_1
X_7611_ _7611_/A _7611_/B VGND VGND VPWR VPWR _7612_/B sky130_fd_sc_hd__nor2_1
X_4823_ _5628_/A VGND VGND VPWR VPWR _5336_/S sky130_fd_sc_hd__buf_2
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4754_ _4817_/S _4757_/B VGND VGND VPWR VPWR _4828_/B sky130_fd_sc_hd__and2_1
X_7542_ _7542_/A _7542_/B VGND VGND VPWR VPWR _7543_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7473_ _7473_/A _7473_/B VGND VGND VPWR VPWR _7474_/C sky130_fd_sc_hd__xnor2_1
X_9212_ _9212_/CLK _9212_/D VGND VGND VPWR VPWR _9212_/Q sky130_fd_sc_hd__dfxtp_2
X_4685_ _4759_/A VGND VGND VPWR VPWR _4966_/B sky130_fd_sc_hd__clkbuf_2
X_6424_ _7037_/A _6907_/A _6607_/A _6424_/D VGND VGND VPWR VPWR _6425_/B sky130_fd_sc_hd__and4_1
X_6355_ _7728_/B VGND VGND VPWR VPWR _7847_/A sky130_fd_sc_hd__buf_2
X_9143_ _9214_/CLK _9143_/D VGND VGND VPWR VPWR _9143_/Q sky130_fd_sc_hd__dfxtp_1
X_9074_ _9214_/CLK _9074_/D VGND VGND VPWR VPWR _9074_/Q sky130_fd_sc_hd__dfxtp_1
X_5306_ _5696_/S VGND VGND VPWR VPWR _5427_/S sky130_fd_sc_hd__clkbuf_2
X_6286_ _6377_/A _6286_/B VGND VGND VPWR VPWR _6288_/A sky130_fd_sc_hd__nor2_1
XFILLER_102_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8025_ _8025_/A _8025_/B VGND VGND VPWR VPWR _9094_/D sky130_fd_sc_hd__xnor2_1
X_5237_ _5122_/X _5236_/X _5305_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5168_ _5132_/X _5532_/A _5163_/X _5167_/Y _4642_/A VGND VGND VPWR VPWR _5168_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5099_ _4535_/A _5096_/X _5097_/Y _5098_/X _5743_/S VGND VGND VPWR VPWR _5099_/X
+ sky130_fd_sc_hd__o221a_1
X_8927_ _9004_/A _8975_/A VGND VGND VPWR VPWR _8929_/C sky130_fd_sc_hd__and2_1
XFILLER_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8858_ _8859_/A _8859_/B VGND VGND VPWR VPWR _8908_/A sky130_fd_sc_hd__nand2_1
X_8789_ _8726_/A _8726_/B _8729_/B VGND VGND VPWR VPWR _8790_/B sky130_fd_sc_hd__a21o_1
X_7809_ _7810_/C _7810_/B _7807_/Y _7808_/X VGND VGND VPWR VPWR _7811_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6140_ _6325_/A _6925_/A _7148_/B _6325_/B VGND VGND VPWR VPWR _6145_/C sky130_fd_sc_hd__a22o_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6071_/A _6071_/B _6071_/C VGND VGND VPWR VPWR _6087_/C sky130_fd_sc_hd__nand3_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _4999_/X _4972_/Y _5019_/X _5021_/X VGND VGND VPWR VPWR _5022_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6973_ _6924_/A _6923_/A _6923_/B VGND VGND VPWR VPWR _7077_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5924_ _7349_/A VGND VGND VPWR VPWR _7131_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8712_ _8770_/B _8771_/A VGND VGND VPWR VPWR _8773_/B sky130_fd_sc_hd__or2_1
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8643_ _8644_/A _8644_/B VGND VGND VPWR VPWR _8645_/A sky130_fd_sc_hd__nand2_1
X_5855_ _5854_/A _5854_/C _5854_/B VGND VGND VPWR VPWR _5858_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4806_ _4891_/A _4836_/A _4980_/A VGND VGND VPWR VPWR _4806_/Y sky130_fd_sc_hd__a21oi_1
X_8574_ _8501_/B _8572_/Y _8570_/Y _8642_/B VGND VGND VPWR VPWR _8648_/A sky130_fd_sc_hd__o211ai_4
X_5786_ _5786_/A VGND VGND VPWR VPWR _9151_/D sky130_fd_sc_hd__buf_4
X_7525_ _7379_/X _7382_/A _7661_/B _7523_/Y VGND VGND VPWR VPWR _7665_/A sky130_fd_sc_hd__a211oi_4
X_4737_ _4737_/A VGND VGND VPWR VPWR _4737_/X sky130_fd_sc_hd__clkbuf_2
X_7456_ _7730_/A VGND VGND VPWR VPWR _8175_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4668_ _9091_/Q VGND VGND VPWR VPWR _5244_/A sky130_fd_sc_hd__clkbuf_2
X_6407_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6409_/A sky130_fd_sc_hd__xnor2_1
X_9126_ _9218_/CLK hold3/X VGND VGND VPWR VPWR _9126_/Q sky130_fd_sc_hd__dfxtp_1
X_4599_ _4599_/A VGND VGND VPWR VPWR _4600_/A sky130_fd_sc_hd__clkbuf_2
X_7387_ _7385_/Y _7386_/X _7277_/D _7277_/Y VGND VGND VPWR VPWR _7539_/B sky130_fd_sc_hd__a211o_1
X_6338_ _6572_/B _6680_/A _6907_/B _7199_/A VGND VGND VPWR VPWR _6340_/A sky130_fd_sc_hd__a22oi_1
X_6269_ _9204_/Q VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9057_ _9057_/A _9057_/B VGND VGND VPWR VPWR _9058_/A sky130_fd_sc_hd__and2_1
X_8008_ _8008_/A _8008_/B VGND VGND VPWR VPWR _8011_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5640_ _5244_/A _4667_/A _5638_/X _5639_/Y _4600_/A VGND VGND VPWR VPWR _5640_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5571_ _4573_/A _4966_/A _5570_/X VGND VGND VPWR VPWR _5571_/Y sky130_fd_sc_hd__o21ai_1
X_8290_ _8290_/A VGND VGND VPWR VPWR _8530_/A sky130_fd_sc_hd__clkbuf_2
X_7310_ _7310_/A _7310_/B VGND VGND VPWR VPWR _7441_/B sky130_fd_sc_hd__xnor2_1
X_7241_ _9201_/Q _7241_/B VGND VGND VPWR VPWR _7245_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7172_ _7172_/A _7172_/B _7172_/C VGND VGND VPWR VPWR _7176_/B sky130_fd_sc_hd__and3_1
X_6123_ _6123_/A _6131_/A VGND VGND VPWR VPWR _6124_/B sky130_fd_sc_hd__nor2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6054_ _6139_/A VGND VGND VPWR VPWR _6223_/A sky130_fd_sc_hd__clkbuf_4
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5146_/A _4937_/A _4933_/A _5656_/B VGND VGND VPWR VPWR _5005_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6956_ _6957_/A _6957_/B VGND VGND VPWR VPWR _6956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5907_ _9168_/Q VGND VGND VPWR VPWR _6702_/A sky130_fd_sc_hd__clkbuf_2
X_6887_ _9180_/Q VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8626_ _8552_/B _8556_/C _8623_/Y _8624_/X VGND VGND VPWR VPWR _8627_/A sky130_fd_sc_hd__a211oi_2
X_5838_ _6235_/A VGND VGND VPWR VPWR _7359_/A sky130_fd_sc_hd__buf_2
X_8557_ _8555_/Y _8635_/A _8478_/B _8480_/X VGND VGND VPWR VPWR _8559_/B sky130_fd_sc_hd__o211a_1
X_5769_ _4635_/A _5768_/Y _4872_/S VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__o21a_1
X_7508_ _9184_/Q VGND VGND VPWR VPWR _7769_/A sky130_fd_sc_hd__clkbuf_2
X_8488_ _8487_/B _8565_/B _8487_/A VGND VGND VPWR VPWR _8489_/B sky130_fd_sc_hd__o21a_1
X_7439_ _7439_/A _7590_/B VGND VGND VPWR VPWR _7440_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9109_ _9218_/CLK _9109_/D VGND VGND VPWR VPWR _9109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6810_ _6810_/A _6810_/B _6810_/C VGND VGND VPWR VPWR _6940_/C sky130_fd_sc_hd__and3_2
X_7790_ _7790_/A _7790_/B VGND VGND VPWR VPWR _7791_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6741_ _6845_/A _6845_/B VGND VGND VPWR VPWR _6743_/A sky130_fd_sc_hd__and2_1
X_6672_ _6597_/A _6596_/B _6596_/A VGND VGND VPWR VPWR _6773_/A sky130_fd_sc_hd__o21ba_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8411_ _8415_/A _9029_/A _8286_/A _8410_/X VGND VGND VPWR VPWR _8411_/Y sky130_fd_sc_hd__a31oi_1
X_5623_ _5749_/A _5403_/X _5620_/X _5622_/Y _4770_/X VGND VGND VPWR VPWR _5623_/X
+ sky130_fd_sc_hd__a221o_1
X_8342_ _8343_/A _8470_/A _8343_/C VGND VGND VPWR VPWR _8344_/A sky130_fd_sc_hd__o21a_1
X_5554_ _5509_/X _5553_/X _5603_/S VGND VGND VPWR VPWR _5554_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8273_ _8792_/D VGND VGND VPWR VPWR _8844_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5485_ _5485_/A _5634_/B VGND VGND VPWR VPWR _5485_/Y sky130_fd_sc_hd__nand2_1
X_7224_ _7224_/A _7224_/B VGND VGND VPWR VPWR _7233_/A sky130_fd_sc_hd__xnor2_1
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7155_ _7230_/B _7155_/B VGND VGND VPWR VPWR _7237_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6036_/C _6036_/Y _6103_/X _6104_/Y VGND VGND VPWR VPWR _6118_/C sky130_fd_sc_hd__o211ai_2
X_7086_ _7086_/A _7205_/B VGND VGND VPWR VPWR _7087_/B sky130_fd_sc_hd__xnor2_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6037_ _6037_/A _6037_/B _6037_/C VGND VGND VPWR VPWR _6037_/Y sky130_fd_sc_hd__nand3_1
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7988_ _7988_/A _7988_/B VGND VGND VPWR VPWR _7990_/C sky130_fd_sc_hd__and2_1
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6939_ _6939_/A _6939_/B _7054_/A VGND VGND VPWR VPWR _6939_/X sky130_fd_sc_hd__or3_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8609_ _8733_/A _8724_/A _8610_/C VGND VGND VPWR VPWR _8661_/B sky130_fd_sc_hd__a21oi_1
XFILLER_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5270_ _5713_/S _5184_/X _5269_/X _5714_/S VGND VGND VPWR VPWR _5270_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8960_ _8859_/A _8859_/B _8908_/B _8959_/Y VGND VGND VPWR VPWR _8973_/B sky130_fd_sc_hd__a31o_1
X_7911_ _7911_/A _7911_/B VGND VGND VPWR VPWR _8018_/B sky130_fd_sc_hd__nand2_1
X_8891_ _8974_/A _8891_/B VGND VGND VPWR VPWR _8925_/A sky130_fd_sc_hd__and2_1
X_7842_ _7842_/A _7915_/B VGND VGND VPWR VPWR _7898_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7773_ _7772_/A _7772_/B _7772_/C VGND VGND VPWR VPWR _7891_/A sky130_fd_sc_hd__o21ai_1
X_4985_ _4985_/A VGND VGND VPWR VPWR _9156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6724_ _6831_/A _6831_/B VGND VGND VPWR VPWR _6730_/B sky130_fd_sc_hd__or2_1
X_6655_ _6655_/A _6655_/B _6655_/C VGND VGND VPWR VPWR _6748_/A sky130_fd_sc_hd__and3_1
X_6586_ _7499_/A _7602_/A VGND VGND VPWR VPWR _6592_/A sky130_fd_sc_hd__nand2_1
X_5606_ _5606_/A VGND VGND VPWR VPWR _5606_/X sky130_fd_sc_hd__clkbuf_2
X_8325_ _8325_/A _8421_/A _8325_/C VGND VGND VPWR VPWR _8325_/X sky130_fd_sc_hd__or3_1
X_5537_ _5149_/A _5210_/A _4586_/A VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8256_ _8256_/A _8398_/B VGND VGND VPWR VPWR _8257_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5468_ _5003_/X _5124_/A _4597_/A VGND VGND VPWR VPWR _5468_/Y sky130_fd_sc_hd__a21oi_1
X_7207_ _7208_/A _7208_/B VGND VGND VPWR VPWR _7209_/A sky130_fd_sc_hd__nand2_1
X_8187_ _8371_/A _8782_/A _8053_/A _8051_/B VGND VGND VPWR VPWR _8196_/A sky130_fd_sc_hd__a31o_1
X_5399_ _5339_/X _5398_/X _5481_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7138_ _7139_/B _7139_/C _7139_/A VGND VGND VPWR VPWR _7140_/A sky130_fd_sc_hd__a21o_1
XFILLER_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7069_ _7064_/A _6957_/X _7064_/B VGND VGND VPWR VPWR _7070_/A sky130_fd_sc_hd__a21boi_1
XFILLER_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 A[26] VGND VGND VPWR VPWR _9188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4770_ _9107_/Q VGND VGND VPWR VPWR _4770_/X sky130_fd_sc_hd__buf_2
X_6440_ _7359_/A VGND VGND VPWR VPWR _7016_/A sky130_fd_sc_hd__clkbuf_2
X_6371_ _6372_/B _6372_/C _6372_/A VGND VGND VPWR VPWR _6375_/A sky130_fd_sc_hd__o21ai_1
X_8110_ _8111_/A _8217_/B _8111_/C VGND VGND VPWR VPWR _8112_/A sky130_fd_sc_hd__o21ai_1
X_5322_ _5158_/A _5555_/A _5320_/X _5321_/Y _5135_/A VGND VGND VPWR VPWR _5322_/X
+ sky130_fd_sc_hd__a221o_1
X_9090_ _9090_/CLK _9090_/D VGND VGND VPWR VPWR _9090_/Q sky130_fd_sc_hd__dfxtp_1
X_8041_ _8041_/A _8041_/B VGND VGND VPWR VPWR _8215_/B sky130_fd_sc_hd__xnor2_1
X_5253_ _5371_/A _5362_/A _4571_/A VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__o21a_1
X_5184_ _5184_/A VGND VGND VPWR VPWR _5184_/X sky130_fd_sc_hd__buf_2
XFILLER_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8943_ _9015_/B _8943_/B VGND VGND VPWR VPWR _8954_/A sky130_fd_sc_hd__or2_1
X_8874_ _8874_/A _8874_/B VGND VGND VPWR VPWR _8876_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7825_ _7935_/C _7825_/B VGND VGND VPWR VPWR _7934_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7756_ _7756_/A VGND VGND VPWR VPWR _8148_/A sky130_fd_sc_hd__clkbuf_2
X_4968_ _4880_/A _4965_/X _4966_/X _4967_/X VGND VGND VPWR VPWR _4968_/Y sky130_fd_sc_hd__o211ai_1
X_7687_ _7686_/A _7686_/B _7685_/Y VGND VGND VPWR VPWR _7688_/B sky130_fd_sc_hd__o21ba_1
X_6707_ _6574_/B _6576_/B _6574_/A VGND VGND VPWR VPWR _6708_/B sky130_fd_sc_hd__o21ba_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4899_ _5676_/B _4882_/B _5337_/B VGND VGND VPWR VPWR _4899_/Y sky130_fd_sc_hd__a21boi_1
X_6638_ _6744_/A _6638_/B VGND VGND VPWR VPWR _6640_/A sky130_fd_sc_hd__and2_1
XFILLER_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8308_ _8306_/X _8307_/Y _8165_/B _8168_/C VGND VGND VPWR VPWR _8308_/X sky130_fd_sc_hd__o211a_1
X_6569_ _6569_/A _6569_/B VGND VGND VPWR VPWR _6571_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8239_ _8517_/A _8337_/A _8542_/C _8239_/D VGND VGND VPWR VPWR _8240_/B sky130_fd_sc_hd__and4_1
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5940_ _5940_/A VGND VGND VPWR VPWR _7093_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7610_ _7852_/A _7610_/B _7610_/C _7610_/D VGND VGND VPWR VPWR _7611_/B sky130_fd_sc_hd__and4_1
XFILLER_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5871_ _5871_/A _5871_/B VGND VGND VPWR VPWR _5881_/A sky130_fd_sc_hd__xnor2_2
X_8590_ _8590_/A _8668_/B VGND VGND VPWR VPWR _8591_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ _5742_/S VGND VGND VPWR VPWR _5628_/A sky130_fd_sc_hd__clkbuf_2
X_4753_ _4842_/B _4753_/B VGND VGND VPWR VPWR _4757_/B sky130_fd_sc_hd__nand2_1
X_7541_ _7539_/C _7539_/Y _7537_/X _7668_/B VGND VGND VPWR VPWR _7542_/B sky130_fd_sc_hd__a211o_1
X_7472_ _7618_/B _7472_/B VGND VGND VPWR VPWR _7473_/B sky130_fd_sc_hd__xnor2_1
X_6423_ _7869_/A _7435_/A _7628_/A _7146_/A VGND VGND VPWR VPWR _6425_/A sky130_fd_sc_hd__a22oi_2
X_4684_ _4688_/A _4688_/B VGND VGND VPWR VPWR _4759_/A sky130_fd_sc_hd__and2_2
X_9211_ _9214_/CLK _9211_/D VGND VGND VPWR VPWR _9211_/Q sky130_fd_sc_hd__dfxtp_2
X_6354_ _7327_/C VGND VGND VPWR VPWR _7728_/B sky130_fd_sc_hd__clkbuf_2
X_9142_ _9219_/CLK _9142_/D VGND VGND VPWR VPWR _9142_/Q sky130_fd_sc_hd__dfxtp_1
X_9073_ _9214_/CLK _9073_/D VGND VGND VPWR VPWR _9073_/Q sky130_fd_sc_hd__dfxtp_2
X_6285_ _6285_/A _6285_/B _6285_/C VGND VGND VPWR VPWR _6286_/B sky130_fd_sc_hd__and3_1
X_5305_ _5120_/X _5304_/X _5305_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8024_ _8024_/A _8024_/B VGND VGND VPWR VPWR _8025_/B sky130_fd_sc_hd__nand2_1
X_5236_ _5208_/X _5235_/X _5236_/S VGND VGND VPWR VPWR _5236_/X sky130_fd_sc_hd__mux2_1
X_5167_ _5165_/X _5166_/Y _4607_/A VGND VGND VPWR VPWR _5167_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5098_ _4980_/B _5028_/A _5043_/A _5742_/S VGND VGND VPWR VPWR _5098_/X sky130_fd_sc_hd__a31o_1
X_8926_ _8978_/A _8926_/B _9002_/A VGND VGND VPWR VPWR _8929_/B sky130_fd_sc_hd__nand3_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8857_ _8790_/A _8790_/B _8804_/B VGND VGND VPWR VPWR _8859_/B sky130_fd_sc_hd__a21bo_1
X_8788_ _8839_/A _8788_/B VGND VGND VPWR VPWR _8790_/A sky130_fd_sc_hd__nor2_1
X_7808_ _7925_/A _7808_/B _7923_/C _7923_/D VGND VGND VPWR VPWR _7808_/X sky130_fd_sc_hd__and4_1
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7739_ _7739_/A _7739_/B VGND VGND VPWR VPWR _7740_/C sky130_fd_sc_hd__xnor2_1
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6071_/A _6071_/B _6071_/C VGND VGND VPWR VPWR _6087_/B sky130_fd_sc_hd__a21o_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5020_/X _4937_/X _5187_/A VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8711_ _8645_/B _8709_/X _8707_/X _8768_/B VGND VGND VPWR VPWR _8771_/A sky130_fd_sc_hd__a211oi_1
X_6972_ _6968_/A _8185_/A _6862_/B _6861_/A VGND VGND VPWR VPWR _7078_/A sky130_fd_sc_hd__a31o_1
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5923_ _9199_/Q VGND VGND VPWR VPWR _7349_/A sky130_fd_sc_hd__clkbuf_2
X_8642_ _8571_/B _8642_/B VGND VGND VPWR VPWR _8644_/B sky130_fd_sc_hd__and2b_1
X_5854_ _5854_/A _5854_/B _5854_/C VGND VGND VPWR VPWR _5858_/A sky130_fd_sc_hd__or3_1
X_8573_ _8570_/Y _8642_/B _8501_/B _8572_/Y VGND VGND VPWR VPWR _8573_/X sky130_fd_sc_hd__a211o_1
X_4805_ _9111_/Q VGND VGND VPWR VPWR _4980_/A sky130_fd_sc_hd__clkbuf_2
X_7524_ _7661_/B _7523_/Y _7379_/X _7382_/A VGND VGND VPWR VPWR _7527_/C sky130_fd_sc_hd__o211a_2
X_5785_ _5117_/X _5784_/X _5785_/S VGND VGND VPWR VPWR _5786_/A sky130_fd_sc_hd__mux2_1
X_4736_ _4769_/A _4736_/B VGND VGND VPWR VPWR _4736_/Y sky130_fd_sc_hd__nor2_1
X_7455_ _7455_/A VGND VGND VPWR VPWR _7730_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4667_ _4667_/A VGND VGND VPWR VPWR _5460_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6406_ _6406_/A _6406_/B VGND VGND VPWR VPWR _6407_/B sky130_fd_sc_hd__nor2_1
X_7386_ _7386_/A _7533_/B _7386_/C VGND VGND VPWR VPWR _7386_/X sky130_fd_sc_hd__or3_4
X_6337_ _7348_/A VGND VGND VPWR VPWR _6680_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9125_ _9220_/CLK hold10/X VGND VGND VPWR VPWR _9125_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4598_ _4598_/A VGND VGND VPWR VPWR _4599_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9056_ _9056_/A _9060_/B VGND VGND VPWR VPWR _9057_/B sky130_fd_sc_hd__or2_1
X_6268_ _6268_/A _6181_/B VGND VGND VPWR VPWR _6285_/B sky130_fd_sc_hd__or2b_1
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8007_ _8007_/A _8007_/B VGND VGND VPWR VPWR _8008_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6199_ _6572_/D VGND VGND VPWR VPWR _7610_/B sky130_fd_sc_hd__buf_2
X_5219_ _5219_/A VGND VGND VPWR VPWR _5219_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8909_ _8909_/A _8909_/B VGND VGND VPWR VPWR _8959_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_clk clkbuf_4_1_0_clk/A VGND VGND VPWR VPWR _9199_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5570_ _5558_/X _4548_/A _5568_/X _5569_/Y _5230_/X VGND VGND VPWR VPWR _5570_/X
+ sky130_fd_sc_hd__a221o_1
X_7240_ _7133_/A _7132_/A _7132_/B VGND VGND VPWR VPWR _7324_/A sky130_fd_sc_hd__o21ba_1
X_7171_ _7171_/A _7171_/B VGND VGND VPWR VPWR _7172_/C sky130_fd_sc_hd__nand2_1
XFILLER_58_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6122_ _6221_/A VGND VGND VPWR VPWR _6123_/A sky130_fd_sc_hd__inv_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6053_ _6053_/A _6053_/B VGND VGND VPWR VPWR _9075_/D sky130_fd_sc_hd__xnor2_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _4940_/A _4842_/A _4783_/A VGND VGND VPWR VPWR _5004_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6955_ _7066_/A _6955_/B VGND VGND VPWR VPWR _9085_/D sky130_fd_sc_hd__xnor2_1
XFILLER_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5906_ _5906_/A _5906_/B _5906_/C VGND VGND VPWR VPWR _5915_/B sky130_fd_sc_hd__nand3_1
X_8625_ _8623_/Y _8624_/X _8552_/B _8556_/C VGND VGND VPWR VPWR _8628_/B sky130_fd_sc_hd__o211ai_2
X_6886_ _6886_/A _6886_/B _7503_/C VGND VGND VPWR VPWR _6891_/B sky130_fd_sc_hd__nand3_1
X_5837_ _6256_/A VGND VGND VPWR VPWR _7083_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8556_ _8556_/A _8556_/B _8556_/C VGND VGND VPWR VPWR _8635_/A sky130_fd_sc_hd__and3_2
X_5768_ _4661_/A _4573_/A _5747_/Y _5450_/A _5432_/A VGND VGND VPWR VPWR _5768_/Y
+ sky130_fd_sc_hd__a221oi_2
X_7507_ _7507_/A _7651_/A VGND VGND VPWR VPWR _7645_/C sky130_fd_sc_hd__nor2_1
X_8487_ _8487_/A _8487_/B _8565_/B VGND VGND VPWR VPWR _8562_/A sky130_fd_sc_hd__nor3_1
X_4719_ _4923_/A _4693_/Y _5071_/A _4721_/A VGND VGND VPWR VPWR _4719_/X sky130_fd_sc_hd__a211o_1
X_7438_ _7438_/A _7438_/B VGND VGND VPWR VPWR _7590_/B sky130_fd_sc_hd__xnor2_1
X_5699_ _5676_/B _5698_/X _5204_/A _4999_/X VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7369_ _7369_/A _7369_/B VGND VGND VPWR VPWR _7495_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9108_ _9218_/CLK _9108_/D VGND VGND VPWR VPWR _9108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9039_ _9022_/A _9022_/B _9038_/Y VGND VGND VPWR VPWR _9040_/B sky130_fd_sc_hd__o21ai_1
XFILLER_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6740_ _6740_/A _6740_/B _6740_/C VGND VGND VPWR VPWR _6845_/B sky130_fd_sc_hd__nand3_2
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6671_ _6671_/A _6671_/B VGND VGND VPWR VPWR _6673_/A sky130_fd_sc_hd__xnor2_1
X_8410_ _8284_/B _8410_/B VGND VGND VPWR VPWR _8410_/X sky130_fd_sc_hd__and2b_1
X_5622_ _5621_/X _5126_/X _5181_/X VGND VGND VPWR VPWR _5622_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8341_ _8584_/A _8733_/A VGND VGND VPWR VPWR _8343_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_5553_ _5484_/X _5552_/X _5553_/S VGND VGND VPWR VPWR _5553_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8272_ _8595_/D VGND VGND VPWR VPWR _8792_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5484_ _5484_/A VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7223_ _7223_/A _7223_/B VGND VGND VPWR VPWR _7224_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _6143_/B _7153_/D _7151_/Y _7230_/A VGND VGND VPWR VPWR _7155_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6103_/X _6104_/Y _6036_/C _6036_/Y VGND VGND VPWR VPWR _6118_/B sky130_fd_sc_hd__a211o_1
X_7085_ _7085_/A _7085_/B VGND VGND VPWR VPWR _7205_/B sky130_fd_sc_hd__xnor2_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A _6036_/B _6036_/C VGND VGND VPWR VPWR _6036_/Y sky130_fd_sc_hd__nor3_2
XFILLER_27_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer20 _5862_/X VGND VGND VPWR VPWR _5931_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7987_ _8068_/A _8257_/C VGND VGND VPWR VPWR _7990_/B sky130_fd_sc_hd__or2_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _6939_/B _7054_/A _6939_/A VGND VGND VPWR VPWR _6938_/Y sky130_fd_sc_hd__o21ai_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6869_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6877_/A sky130_fd_sc_hd__nand2_1
X_8608_ _8608_/A _8662_/A VGND VGND VPWR VPWR _8610_/C sky130_fd_sc_hd__nor2_1
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8539_ _8816_/A _8832_/A _8469_/A _8465_/B VGND VGND VPWR VPWR _8548_/A sky130_fd_sc_hd__a31o_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8890_ _8890_/A _8890_/B VGND VGND VPWR VPWR _8902_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7910_ _8022_/A _7910_/B VGND VGND VPWR VPWR _9093_/D sky130_fd_sc_hd__xnor2_1
X_7841_ _7841_/A _7841_/B _7841_/C VGND VGND VPWR VPWR _7915_/B sky130_fd_sc_hd__and3_1
XFILLER_91_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7772_ _7772_/A _7772_/B _7772_/C VGND VGND VPWR VPWR _7774_/A sky130_fd_sc_hd__or3_1
XFILLER_63_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4984_ _4971_/B _4983_/X _5653_/B VGND VGND VPWR VPWR _4985_/A sky130_fd_sc_hd__mux2_1
X_6723_ _7093_/B _7583_/D VGND VGND VPWR VPWR _6831_/B sky130_fd_sc_hd__nand2_2
X_6654_ _6654_/A _6654_/B VGND VGND VPWR VPWR _6747_/A sky130_fd_sc_hd__and2_1
X_5605_ _5583_/X _5510_/X _5511_/X _5603_/X _5604_/X VGND VGND VPWR VPWR _9143_/D
+ sky130_fd_sc_hd__o221a_2
X_6585_ _6585_/A _6585_/B VGND VGND VPWR VPWR _6601_/B sky130_fd_sc_hd__nand2_1
X_8324_ _8325_/A _8421_/A _8325_/C VGND VGND VPWR VPWR _8324_/Y sky130_fd_sc_hd__o21ai_1
X_5536_ _5179_/A _5369_/A _5535_/X VGND VGND VPWR VPWR _5536_/Y sky130_fd_sc_hd__a21oi_1
X_8255_ _8255_/A _8255_/B VGND VGND VPWR VPWR _8398_/B sky130_fd_sc_hd__nor2_1
X_5467_ _5215_/X _5184_/A _5465_/X _5466_/Y _5222_/X VGND VGND VPWR VPWR _5467_/X
+ sky130_fd_sc_hd__a221o_1
X_7206_ _7087_/A _7087_/B _7205_/X VGND VGND VPWR VPWR _7208_/B sky130_fd_sc_hd__a21oi_1
X_8186_ _8724_/A VGND VGND VPWR VPWR _8782_/A sky130_fd_sc_hd__clkbuf_4
X_5398_ _5315_/X _5397_/X _5428_/S VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7137_ _7219_/A _7137_/B VGND VGND VPWR VPWR _7139_/A sky130_fd_sc_hd__xnor2_2
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7068_ _7068_/A _7068_/B VGND VGND VPWR VPWR _7071_/B sky130_fd_sc_hd__or2_1
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6019_ _5976_/B _5976_/C _5976_/A VGND VGND VPWR VPWR _6021_/C sky130_fd_sc_hd__a21bo_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6370_ _6370_/A _6370_/B VGND VGND VPWR VPWR _6372_/A sky130_fd_sc_hd__xnor2_1
X_5321_ _4841_/A _5248_/Y _5222_/X VGND VGND VPWR VPWR _5321_/Y sky130_fd_sc_hd__a21oi_1
X_8040_ _8322_/A _8597_/B VGND VGND VPWR VPWR _8041_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5252_ _5252_/A VGND VGND VPWR VPWR _5371_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5183_ _9083_/Q VGND VGND VPWR VPWR _5184_/A sky130_fd_sc_hd__inv_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8942_ _8941_/B _8942_/B VGND VGND VPWR VPWR _8943_/B sky130_fd_sc_hd__and2b_1
XFILLER_71_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8873_ _8872_/A _8872_/B _8872_/C VGND VGND VPWR VPWR _8874_/B sky130_fd_sc_hd__a21oi_1
X_7824_ _7923_/B _7824_/B VGND VGND VPWR VPWR _7825_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7755_ _7629_/B _7752_/Y _7754_/Y VGND VGND VPWR VPWR _7759_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4967_ _4726_/X _5080_/A _4963_/B _5692_/S VGND VGND VPWR VPWR _4967_/X sky130_fd_sc_hd__o31a_1
X_7686_ _7686_/A _7686_/B _7685_/Y VGND VGND VPWR VPWR _7688_/A sky130_fd_sc_hd__nor3b_1
X_6706_ _6706_/A _6706_/B VGND VGND VPWR VPWR _6769_/B sky130_fd_sc_hd__xnor2_1
X_4898_ _5506_/A VGND VGND VPWR VPWR _5337_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6637_ _6637_/A _6637_/B _6637_/C VGND VGND VPWR VPWR _6638_/B sky130_fd_sc_hd__nand3_1
X_6568_ _7421_/C _7847_/A _7459_/D _6700_/A VGND VGND VPWR VPWR _6569_/B sky130_fd_sc_hd__a22oi_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8307_ _8307_/A _8307_/B VGND VGND VPWR VPWR _8307_/Y sky130_fd_sc_hd__nor2_2
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5519_ _5214_/X _5194_/X _5517_/X _5518_/Y _5001_/A VGND VGND VPWR VPWR _5519_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6499_ _6499_/A _6499_/B VGND VGND VPWR VPWR _6507_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8238_ _8337_/A _8542_/C _8239_/D _8587_/A VGND VGND VPWR VPWR _8240_/A sky130_fd_sc_hd__a22oi_1
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8169_ _8168_/B _8168_/C _8168_/A VGND VGND VPWR VPWR _8169_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5870_ _5825_/X _5870_/B VGND VGND VPWR VPWR _5871_/B sky130_fd_sc_hd__and2b_1
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4821_ _9111_/Q VGND VGND VPWR VPWR _5742_/S sky130_fd_sc_hd__inv_2
XFILLER_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4752_ _4842_/B _4753_/B VGND VGND VPWR VPWR _4817_/S sky130_fd_sc_hd__or2_2
X_7540_ _7537_/X _7668_/B _7539_/C _7539_/Y VGND VGND VPWR VPWR _7542_/A sky130_fd_sc_hd__o211ai_1
X_7471_ _7334_/A _7333_/A _7333_/B VGND VGND VPWR VPWR _7472_/B sky130_fd_sc_hd__o21ba_1
X_4683_ _9121_/Q _9113_/Q _4691_/B VGND VGND VPWR VPWR _4688_/B sky130_fd_sc_hd__or3_1
X_9210_ _9210_/CLK _9210_/D VGND VGND VPWR VPWR _9210_/Q sky130_fd_sc_hd__dfxtp_2
X_6422_ _6907_/B VGND VGND VPWR VPWR _7628_/A sky130_fd_sc_hd__buf_2
X_9141_ _9208_/CLK _9141_/D VGND VGND VPWR VPWR _9141_/Q sky130_fd_sc_hd__dfxtp_1
X_6353_ _9205_/Q VGND VGND VPWR VPWR _7327_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9072_ _9090_/CLK _9072_/D VGND VGND VPWR VPWR _9072_/Q sky130_fd_sc_hd__dfxtp_1
X_5304_ _5206_/X _5302_/X _5527_/S VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__mux2_1
X_6284_ _6285_/A _6285_/B _6285_/C VGND VGND VPWR VPWR _6377_/A sky130_fd_sc_hd__a21oi_4
XFILLER_102_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5235_ _5124_/X _5234_/X _5354_/S VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__mux2_1
X_8023_ _7796_/A _7796_/B _7792_/Y _7794_/B _8022_/Y VGND VGND VPWR VPWR _8024_/B
+ sky130_fd_sc_hd__o311ai_4
XFILLER_102_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5166_ _9077_/Q VGND VGND VPWR VPWR _5166_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5097_ _4980_/B _5028_/A _5043_/A VGND VGND VPWR VPWR _5097_/Y sky130_fd_sc_hd__a21oi_1
X_8925_ _8925_/A VGND VGND VPWR VPWR _9002_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8856_ _8856_/A _8904_/B VGND VGND VPWR VPWR _8859_/A sky130_fd_sc_hd__and2_1
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8787_ _8787_/A _8787_/B _8787_/C VGND VGND VPWR VPWR _8788_/B sky130_fd_sc_hd__nor3_1
X_7807_ _7810_/D VGND VGND VPWR VPWR _7807_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5999_ _5999_/A _5999_/B VGND VGND VPWR VPWR _6047_/B sky130_fd_sc_hd__nand2_2
X_7738_ _7843_/B _7738_/B VGND VGND VPWR VPWR _7739_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7669_ _7668_/A _7668_/B _7668_/C VGND VGND VPWR VPWR _7793_/A sky130_fd_sc_hd__o21ai_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5391_/A VGND VGND VPWR VPWR _5020_/X sky130_fd_sc_hd__clkbuf_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6971_ _7940_/B VGND VGND VPWR VPWR _8185_/A sky130_fd_sc_hd__buf_2
XFILLER_65_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8710_ _8707_/X _8768_/B _8645_/B _8709_/X VGND VGND VPWR VPWR _8770_/B sky130_fd_sc_hd__o211a_1
XFILLER_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5922_ _5922_/A VGND VGND VPWR VPWR _7096_/A sky130_fd_sc_hd__clkbuf_2
X_8641_ _8656_/A _8641_/B VGND VGND VPWR VPWR _8644_/A sky130_fd_sc_hd__xor2_1
X_5853_ _6014_/A _7259_/B _6022_/A _6139_/A VGND VGND VPWR VPWR _5854_/C sky130_fd_sc_hd__a22oi_2
X_8572_ _8572_/A VGND VGND VPWR VPWR _8572_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5784_ _4891_/X _4896_/A _5775_/X _5783_/X _4687_/X VGND VGND VPWR VPWR _5784_/X
+ sky130_fd_sc_hd__o32a_1
X_4804_ _4737_/X _4787_/B _4803_/Y _4739_/X VGND VGND VPWR VPWR _4804_/X sky130_fd_sc_hd__a211o_1
X_7523_ _7522_/A _7522_/B _7522_/C VGND VGND VPWR VPWR _7523_/Y sky130_fd_sc_hd__a21oi_2
X_4735_ _4693_/Y _4732_/X _5236_/S VGND VGND VPWR VPWR _4736_/B sky130_fd_sc_hd__mux2_1
X_7454_ _7923_/B _7962_/B VGND VGND VPWR VPWR _7461_/A sky130_fd_sc_hd__nand2_1
X_4666_ _5160_/A VGND VGND VPWR VPWR _4667_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6405_ _7293_/A _6405_/B _6759_/C _6572_/D VGND VGND VPWR VPWR _6406_/B sky130_fd_sc_hd__and4_1
X_7385_ _7386_/A _7533_/B _7386_/C VGND VGND VPWR VPWR _7385_/Y sky130_fd_sc_hd__o21ai_2
X_4597_ _4597_/A VGND VGND VPWR VPWR _4598_/A sky130_fd_sc_hd__clkbuf_2
X_9124_ _9219_/CLK hold11/X VGND VGND VPWR VPWR _9124_/Q sky130_fd_sc_hd__dfxtp_1
X_6336_ _7201_/A _6607_/B VGND VGND VPWR VPWR _6341_/A sky130_fd_sc_hd__nand2_1
X_9055_ _9055_/A _9055_/B VGND VGND VPWR VPWR _9072_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6267_ _6267_/A _6180_/B VGND VGND VPWR VPWR _6285_/A sky130_fd_sc_hd__or2b_1
XFILLER_88_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8006_ _8007_/A _8007_/B VGND VGND VPWR VPWR _8008_/A sky130_fd_sc_hd__and2_1
X_6198_ _7152_/C VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__clkbuf_2
X_5218_ _4847_/A _5362_/A _5217_/X _4584_/A VGND VGND VPWR VPWR _5218_/Y sky130_fd_sc_hd__a211oi_1
X_5149_ _5149_/A VGND VGND VPWR VPWR _5149_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8908_ _8908_/A _8908_/B VGND VGND VPWR VPWR _8959_/A sky130_fd_sc_hd__xor2_2
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8839_ _8839_/A _8839_/B VGND VGND VPWR VPWR _8904_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7170_ _7170_/A _7281_/C _7167_/X _7168_/Y VGND VGND VPWR VPWR _7171_/B sky130_fd_sc_hd__or4bb_1
X_6121_ _6213_/A _6213_/B VGND VGND VPWR VPWR _6221_/B sky130_fd_sc_hd__xnor2_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6052_ _9052_/B _9052_/C VGND VGND VPWR VPWR _6053_/B sky130_fd_sc_hd__or2_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5058_/A VGND VGND VPWR VPWR _5003_/X sky130_fd_sc_hd__clkbuf_2
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6954_ _6747_/A _6952_/X _7068_/A VGND VGND VPWR VPWR _6955_/B sky130_fd_sc_hd__o21ai_1
X_5905_ _5906_/A _5906_/B _5906_/C VGND VGND VPWR VPWR _5915_/A sky130_fd_sc_hd__a21o_1
X_8624_ _8624_/A _8624_/B _8624_/C VGND VGND VPWR VPWR _8624_/X sky130_fd_sc_hd__and3_1
X_6885_ _6885_/A _9180_/Q VGND VGND VPWR VPWR _7503_/C sky130_fd_sc_hd__and2_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5836_ _9167_/Q VGND VGND VPWR VPWR _6256_/A sky130_fd_sc_hd__clkbuf_2
X_8555_ _8556_/B _8556_/C _8556_/A VGND VGND VPWR VPWR _8555_/Y sky130_fd_sc_hd__a21oi_2
X_5767_ _5120_/X _4812_/X _5204_/A _5761_/X _5766_/X VGND VGND VPWR VPWR _9150_/D
+ sky130_fd_sc_hd__o221a_1
X_7506_ _7506_/A _7506_/B _7640_/A _7986_/B VGND VGND VPWR VPWR _7651_/A sky130_fd_sc_hd__and4_1
X_8486_ _8395_/B _8397_/X _8483_/Y _8565_/A VGND VGND VPWR VPWR _8565_/B sky130_fd_sc_hd__a211oi_4
X_4718_ _4774_/A VGND VGND VPWR VPWR _4923_/A sky130_fd_sc_hd__clkbuf_2
X_5698_ _5765_/A _5697_/X _5698_/S VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__mux2_1
X_7437_ _7810_/C _7940_/B VGND VGND VPWR VPWR _7438_/B sky130_fd_sc_hd__nand2_1
X_4649_ _5149_/A VGND VGND VPWR VPWR _4650_/A sky130_fd_sc_hd__buf_2
X_7368_ _7368_/A _7368_/B VGND VGND VPWR VPWR _7369_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6319_ _7766_/A _7808_/B _8050_/A _5945_/A VGND VGND VPWR VPWR _6320_/B sky130_fd_sc_hd__a22oi_2
X_9107_ _9219_/CLK _9107_/D VGND VGND VPWR VPWR _9107_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7299_ _7299_/A _9214_/Q VGND VGND VPWR VPWR _7301_/B sky130_fd_sc_hd__and2_1
X_9038_ _9038_/A _9038_/B VGND VGND VPWR VPWR _9038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6670_ _6670_/A _6670_/B VGND VGND VPWR VPWR _6671_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5621_ _5621_/A VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__buf_2
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8340_ _8587_/A _8438_/B _8717_/A _8664_/C VGND VGND VPWR VPWR _8470_/A sky130_fd_sc_hd__and4_1
X_5552_ _5461_/X _5551_/X _5552_/S VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__mux2_1
X_8271_ _8450_/C VGND VGND VPWR VPWR _8978_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5483_ _5461_/X _5365_/X _5366_/X _5481_/X _5482_/X VGND VGND VPWR VPWR _9138_/D
+ sky130_fd_sc_hd__o221a_1
X_7222_ _7325_/A _7453_/A _7222_/C _7222_/D VGND VGND VPWR VPWR _7223_/B sky130_fd_sc_hd__and4_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7153_ _7151_/Y _7230_/A _7153_/C _7153_/D VGND VGND VPWR VPWR _7230_/B sky130_fd_sc_hd__and4bb_1
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7084_ _7084_/A _7084_/B VGND VGND VPWR VPWR _7085_/B sky130_fd_sc_hd__nor2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6104_/A _6104_/B _6104_/C VGND VGND VPWR VPWR _6104_/Y sky130_fd_sc_hd__nand3_2
XFILLER_100_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6036_/B _6036_/C _6036_/A VGND VGND VPWR VPWR _6035_/X sky130_fd_sc_hd__o21a_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer21 _5931_/A1 VGND VGND VPWR VPWR _5932_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7986_ _7986_/A _7986_/B VGND VGND VPWR VPWR _8257_/C sky130_fd_sc_hd__nand2_2
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _6961_/A _6961_/B VGND VGND VPWR VPWR _6939_/A sky130_fd_sc_hd__xnor2_1
X_6868_ _6868_/A _6868_/B VGND VGND VPWR VPWR _6869_/B sky130_fd_sc_hd__or2_1
X_8607_ _8721_/A _8607_/B _8607_/C _8607_/D VGND VGND VPWR VPWR _8662_/A sky130_fd_sc_hd__and4_1
X_5819_ _9162_/Q VGND VGND VPWR VPWR _6031_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8538_ _8538_/A VGND VGND VPWR VPWR _8816_/A sky130_fd_sc_hd__clkbuf_2
X_6799_ _7348_/A _7019_/B _7152_/B _7152_/D VGND VGND VPWR VPWR _6801_/A sky130_fd_sc_hd__and4_1
XFILLER_10_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8469_ _8469_/A _8469_/B VGND VGND VPWR VPWR _8470_/C sky130_fd_sc_hd__xnor2_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput90 _9132_/Q VGND VGND VPWR VPWR F[3] sky130_fd_sc_hd__buf_2
XFILLER_83_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7840_ _7841_/B _7841_/C _7841_/A VGND VGND VPWR VPWR _7842_/A sky130_fd_sc_hd__a21oi_1
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7771_ _7771_/A _7771_/B VGND VGND VPWR VPWR _7772_/C sky130_fd_sc_hd__xnor2_1
X_4983_ _4916_/X _4981_/X _5743_/S VGND VGND VPWR VPWR _4983_/X sky130_fd_sc_hd__mux2_1
X_6722_ _7307_/D VGND VGND VPWR VPWR _7583_/D sky130_fd_sc_hd__clkbuf_2
X_6653_ _6653_/A _6655_/C VGND VGND VPWR VPWR _6654_/A sky130_fd_sc_hd__nand2_1
X_5604_ _5604_/A _5604_/B VGND VGND VPWR VPWR _5604_/X sky130_fd_sc_hd__or2_1
X_6584_ _6584_/A _6539_/A VGND VGND VPWR VPWR _6601_/A sky130_fd_sc_hd__or2b_1
X_8323_ _8323_/A _8423_/B VGND VGND VPWR VPWR _8325_/C sky130_fd_sc_hd__or2_1
X_5535_ _5313_/A _5212_/A _5146_/X _5246_/Y _4856_/A VGND VGND VPWR VPWR _5535_/X
+ sky130_fd_sc_hd__a221o_1
X_8254_ _8254_/A _8254_/B VGND VGND VPWR VPWR _8255_/B sky130_fd_sc_hd__nor2_2
X_5466_ _4862_/A _5211_/A _4591_/A VGND VGND VPWR VPWR _5466_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7205_ _7086_/A _7205_/B VGND VGND VPWR VPWR _7205_/X sky130_fd_sc_hd__and2b_1
X_8185_ _8185_/A VGND VGND VPWR VPWR _8724_/A sky130_fd_sc_hd__buf_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5397_ _5287_/X _5396_/X _5427_/S VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7136_ _7136_/A _7235_/A VGND VGND VPWR VPWR _7137_/B sky130_fd_sc_hd__and2_1
X_7067_ _6654_/A _6654_/B _6952_/X _7068_/B VGND VGND VPWR VPWR _7071_/A sky130_fd_sc_hd__a211o_1
XFILLER_100_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6018_ _6018_/A _6018_/B _6018_/C VGND VGND VPWR VPWR _6021_/B sky130_fd_sc_hd__nand3_1
XFILLER_27_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _8351_/C _8150_/C VGND VGND VPWR VPWR _7970_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A VGND VGND VPWR VPWR clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5320_ _5154_/A _5507_/A _5318_/X _5319_/Y _4591_/A VGND VGND VPWR VPWR _5320_/X
+ sky130_fd_sc_hd__a221o_1
X_5251_ _5251_/A VGND VGND VPWR VPWR _5618_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5182_ _5126_/X _5630_/A _5176_/X _5180_/Y _5181_/X VGND VGND VPWR VPWR _5182_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8941_ _8942_/B _8941_/B VGND VGND VPWR VPWR _9015_/B sky130_fd_sc_hd__and2b_1
XFILLER_56_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8872_ _8872_/A _8872_/B _8872_/C VGND VGND VPWR VPWR _8874_/A sky130_fd_sc_hd__and3_1
X_7823_ _7823_/A _7944_/A VGND VGND VPWR VPWR _7935_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7754_ _7754_/A _7754_/B VGND VGND VPWR VPWR _7754_/Y sky130_fd_sc_hd__nor2_1
X_6705_ _6754_/B _7153_/D VGND VGND VPWR VPWR _6706_/B sky130_fd_sc_hd__nand2_1
X_4966_ _4966_/A _4966_/B _4960_/X VGND VGND VPWR VPWR _4966_/X sky130_fd_sc_hd__or3b_1
X_7685_ _7573_/A _7573_/B _7577_/B VGND VGND VPWR VPWR _7685_/Y sky130_fd_sc_hd__a21oi_1
X_4897_ _4897_/A VGND VGND VPWR VPWR _5506_/A sky130_fd_sc_hd__buf_2
X_6636_ _6637_/A _6637_/B _6637_/C VGND VGND VPWR VPWR _6744_/A sky130_fd_sc_hd__a21o_1
X_6567_ _7187_/A _6567_/B _7604_/C _7847_/C VGND VGND VPWR VPWR _6569_/A sky130_fd_sc_hd__and4_1
X_8306_ _8307_/A _8307_/B VGND VGND VPWR VPWR _8306_/X sky130_fd_sc_hd__and2_1
X_5518_ _5003_/X _5122_/A _4597_/A VGND VGND VPWR VPWR _5518_/Y sky130_fd_sc_hd__a21oi_1
X_6498_ _6968_/B _7962_/B VGND VGND VPWR VPWR _6499_/B sky130_fd_sc_hd__nand2_1
X_8237_ _8162_/A _8162_/B _8236_/X VGND VGND VPWR VPWR _8256_/A sky130_fd_sc_hd__a21oi_1
X_5449_ _5449_/A VGND VGND VPWR VPWR _5450_/A sky130_fd_sc_hd__buf_2
X_8168_ _8168_/A _8168_/B _8168_/C VGND VGND VPWR VPWR _8266_/A sky130_fd_sc_hd__and3_1
X_7119_ _7259_/A _7119_/B _7119_/C _7119_/D VGND VGND VPWR VPWR _7121_/A sky130_fd_sc_hd__and4_1
XFILLER_59_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8099_ _8099_/A _8166_/B VGND VGND VPWR VPWR _8100_/C sky130_fd_sc_hd__or2_1
XFILLER_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4820_ _4914_/A VGND VGND VPWR VPWR _4960_/B sky130_fd_sc_hd__buf_2
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4751_ _9122_/Q _9114_/Q _4688_/A VGND VGND VPWR VPWR _4753_/B sky130_fd_sc_hd__a21boi_1
XFILLER_14_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7470_ _7470_/A _7470_/B VGND VGND VPWR VPWR _7618_/B sky130_fd_sc_hd__xnor2_1
X_4682_ _9121_/Q _9113_/Q _4691_/B VGND VGND VPWR VPWR _4688_/A sky130_fd_sc_hd__o21ai_1
X_6421_ _6321_/A _6320_/B _6320_/A VGND VGND VPWR VPWR _6488_/A sky130_fd_sc_hd__o21ba_2
X_9140_ _9212_/CLK _9140_/D VGND VGND VPWR VPWR _9140_/Q sky130_fd_sc_hd__dfxtp_1
X_6352_ _6261_/A _6352_/B VGND VGND VPWR VPWR _6367_/B sky130_fd_sc_hd__and2b_1
X_9071_ _9090_/CLK _9071_/D VGND VGND VPWR VPWR _9071_/Q sky130_fd_sc_hd__dfxtp_2
X_5303_ _5738_/S VGND VGND VPWR VPWR _5527_/S sky130_fd_sc_hd__clkbuf_2
X_6283_ _6370_/A _6283_/B VGND VGND VPWR VPWR _6285_/C sky130_fd_sc_hd__or2_1
X_8022_ _8022_/A VGND VGND VPWR VPWR _8022_/Y sky130_fd_sc_hd__inv_2
X_5234_ _5653_/A _5232_/Y _5572_/S VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__mux2_1
X_5165_ _5367_/A VGND VGND VPWR VPWR _5165_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5096_ _4739_/X _5092_/X _5094_/Y _5095_/X VGND VGND VPWR VPWR _5096_/X sky130_fd_sc_hd__o22a_1
X_8924_ _8978_/A _8926_/B _8925_/A VGND VGND VPWR VPWR _8929_/A sky130_fd_sc_hd__a21o_1
XFILLER_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8855_ _8855_/A _8855_/B VGND VGND VPWR VPWR _8904_/B sky130_fd_sc_hd__or2_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7806_ _7583_/A _7694_/C _7694_/D _7435_/A VGND VGND VPWR VPWR _7810_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8786_ _8787_/A _8787_/B _8787_/C VGND VGND VPWR VPWR _8839_/A sky130_fd_sc_hd__o21a_1
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5998_ _5997_/B _5997_/C _5997_/A VGND VGND VPWR VPWR _5999_/B sky130_fd_sc_hd__a21o_1
X_7737_ _7612_/A _7611_/A _7611_/B VGND VGND VPWR VPWR _7738_/B sky130_fd_sc_hd__o21ba_1
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4949_ _5621_/A _4946_/X _4948_/Y VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__a21oi_1
X_7668_ _7668_/A _7668_/B _7668_/C VGND VGND VPWR VPWR _7670_/A sky130_fd_sc_hd__or3_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6619_ _6716_/B _6716_/C _6716_/A VGND VGND VPWR VPWR _6619_/Y sky130_fd_sc_hd__o21ai_2
X_7599_ _7684_/A _7599_/B VGND VGND VPWR VPWR _7691_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6970_ _7309_/B VGND VGND VPWR VPWR _7940_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5921_ _7767_/A _6828_/A _5847_/A _5844_/B VGND VGND VPWR VPWR _5961_/C sky130_fd_sc_hd__a31o_1
XFILLER_80_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8640_ _8640_/A _8640_/B VGND VGND VPWR VPWR _8641_/B sky130_fd_sc_hd__and2_1
XFILLER_61_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5852_ _6667_/A VGND VGND VPWR VPWR _7259_/B sky130_fd_sc_hd__clkbuf_4
X_8571_ _8571_/A _8571_/B _8571_/C VGND VGND VPWR VPWR _8642_/B sky130_fd_sc_hd__or3_2
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5783_ _4538_/A _5782_/X _4982_/A VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__o21a_1
X_4803_ _4769_/Y _4802_/X _4737_/A VGND VGND VPWR VPWR _4803_/Y sky130_fd_sc_hd__a21oi_1
X_7522_ _7522_/A _7522_/B _7522_/C VGND VGND VPWR VPWR _7661_/B sky130_fd_sc_hd__and3_2
X_4734_ _5738_/S VGND VGND VPWR VPWR _5236_/S sky130_fd_sc_hd__buf_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7453_ _7453_/A VGND VGND VPWR VPWR _7923_/B sky130_fd_sc_hd__clkbuf_2
X_4665_ _5158_/A VGND VGND VPWR VPWR _5160_/A sky130_fd_sc_hd__clkbuf_2
X_7384_ _7528_/A _7384_/B VGND VGND VPWR VPWR _7386_/C sky130_fd_sc_hd__xor2_2
X_6404_ _7419_/A _6927_/C _6361_/D _6251_/A VGND VGND VPWR VPWR _6406_/A sky130_fd_sc_hd__a22oi_2
X_4596_ _5002_/A VGND VGND VPWR VPWR _4597_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9123_ _9218_/CLK hold17/X VGND VGND VPWR VPWR _9123_/Q sky130_fd_sc_hd__dfxtp_1
X_6335_ _6335_/A _6335_/B VGND VGND VPWR VPWR _6342_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9054_ _9057_/A _9054_/B VGND VGND VPWR VPWR _9055_/B sky130_fd_sc_hd__and2_1
X_8005_ _8005_/A _8005_/B VGND VGND VPWR VPWR _8007_/B sky130_fd_sc_hd__xnor2_1
X_6266_ _6264_/C _6264_/Y _6262_/Y _6263_/X VGND VGND VPWR VPWR _6288_/C sky130_fd_sc_hd__a211o_1
X_6197_ _8091_/A VGND VGND VPWR VPWR _8156_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5217_ _9070_/Q _4579_/A _4659_/A _9069_/Q _5216_/Y VGND VGND VPWR VPWR _5217_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5148_ _5313_/A _9070_/Q _5369_/A _9069_/Q _5147_/X VGND VGND VPWR VPWR _5148_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5079_ _5080_/A _5080_/C _5080_/B VGND VGND VPWR VPWR _5079_/Y sky130_fd_sc_hd__o21ai_1
X_8907_ _8907_/A _8907_/B VGND VGND VPWR VPWR _8908_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8838_ _8839_/A _8839_/B VGND VGND VPWR VPWR _8840_/A sky130_fd_sc_hd__or2_1
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8769_ _8769_/A _8768_/X VGND VGND VPWR VPWR _8880_/A sky130_fd_sc_hd__or2b_1
XFILLER_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6120_ _6041_/A _6041_/B _6041_/C VGND VGND VPWR VPWR _6213_/B sky130_fd_sc_hd__a21bo_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6051_ _6051_/A _6051_/B VGND VGND VPWR VPWR _6053_/A sky130_fd_sc_hd__nor2_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6953_ _6848_/A _6748_/Y _6848_/B VGND VGND VPWR VPWR _7068_/A sky130_fd_sc_hd__a21o_1
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6884_ _6884_/A _6884_/B VGND VGND VPWR VPWR _6901_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5904_ _5854_/B _5854_/C _5854_/A VGND VGND VPWR VPWR _5906_/C sky130_fd_sc_hd__o21bai_1
X_8623_ _8624_/B _8624_/C _8624_/A VGND VGND VPWR VPWR _8623_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5883_/A _5883_/B VGND VGND VPWR VPWR _5863_/C sky130_fd_sc_hd__and2_1
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8554_ _8554_/A _8554_/B VGND VGND VPWR VPWR _8556_/C sky130_fd_sc_hd__or2_2
X_5766_ _5365_/A _5764_/X _5765_/X _4891_/X VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__a31o_1
X_7505_ _6223_/A _7640_/A _7986_/B _6223_/B VGND VGND VPWR VPWR _7507_/A sky130_fd_sc_hd__a22oi_1
X_8485_ _8483_/Y _8565_/A _8395_/B _8397_/X VGND VGND VPWR VPWR _8487_/B sky130_fd_sc_hd__o211a_1
X_5697_ _5632_/X _5696_/X _5697_/S VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__mux2_1
X_4717_ _4714_/X _4698_/X _4717_/S VGND VGND VPWR VPWR _4717_/X sky130_fd_sc_hd__mux2_1
X_7436_ _7436_/A _7436_/B VGND VGND VPWR VPWR _7438_/A sky130_fd_sc_hd__nor2_1
X_4648_ _4856_/A VGND VGND VPWR VPWR _5149_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7367_ _7367_/A _7367_/B _9181_/Q _9182_/Q VGND VGND VPWR VPWR _7368_/B sky130_fd_sc_hd__and4_1
XFILLER_89_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9106_ _9221_/CLK _9106_/D VGND VGND VPWR VPWR _9106_/Q sky130_fd_sc_hd__dfxtp_1
X_4579_ _4579_/A VGND VGND VPWR VPWR _5559_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6318_ _7938_/B VGND VGND VPWR VPWR _8050_/A sky130_fd_sc_hd__buf_2
X_7298_ _7298_/A _7298_/B VGND VGND VPWR VPWR _7301_/A sky130_fd_sc_hd__xor2_1
X_9037_ _9037_/A _9036_/X VGND VGND VPWR VPWR _9040_/A sky130_fd_sc_hd__or2b_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ _6175_/B _6179_/B _6175_/A VGND VGND VPWR VPWR _6261_/A sky130_fd_sc_hd__o21ba_1
XFILLER_103_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5620_ _5402_/A _4656_/A _5617_/X _5619_/Y _5126_/A VGND VGND VPWR VPWR _5620_/X
+ sky130_fd_sc_hd__a221o_1
X_5551_ _5433_/A _4769_/A _5549_/X _5550_/Y VGND VGND VPWR VPWR _5551_/X sky130_fd_sc_hd__a22o_1
X_8270_ _8792_/B VGND VGND VPWR VPWR _8450_/C sky130_fd_sc_hd__clkbuf_1
X_7221_ _7583_/B _6493_/C _7604_/D _7583_/A VGND VGND VPWR VPWR _7223_/A sky130_fd_sc_hd__a22oi_1
X_5482_ _5482_/A _5482_/B VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__or2_1
X_7152_ _7152_/A _7152_/B _7152_/C _7152_/D VGND VGND VPWR VPWR _7230_/A sky130_fd_sc_hd__and4_1
X_7083_ _7083_/A _7083_/B _9208_/Q _7307_/D VGND VGND VPWR VPWR _7084_/B sky130_fd_sc_hd__and4_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6104_/B _6104_/C _6104_/A VGND VGND VPWR VPWR _6103_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6108_/A _6108_/B VGND VGND VPWR VPWR _6036_/A sky130_fd_sc_hd__xnor2_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7985_ _7628_/A _8154_/B _8243_/B _7627_/A VGND VGND VPWR VPWR _7990_/A sky130_fd_sc_hd__a22o_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6936_ _6936_/A _6988_/A VGND VGND VPWR VPWR _6961_/B sky130_fd_sc_hd__nand2_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6867_ _6868_/A _6868_/B VGND VGND VPWR VPWR _6869_/A sky130_fd_sc_hd__nand2_1
X_8606_ _8542_/B _8607_/C _8607_/D _8721_/A VGND VGND VPWR VPWR _8608_/A sky130_fd_sc_hd__a22oi_1
X_6798_ _7129_/A _7153_/C VGND VGND VPWR VPWR _6802_/A sky130_fd_sc_hd__nand2_1
X_5818_ _6055_/A VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__buf_2
XFILLER_10_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8537_ _8537_/A _8537_/B VGND VGND VPWR VPWR _8554_/A sky130_fd_sc_hd__xor2_2
X_5749_ _5749_/A _5749_/B VGND VGND VPWR VPWR _5749_/Y sky130_fd_sc_hd__nor2_1
X_8468_ _8538_/A _8666_/A VGND VGND VPWR VPWR _8469_/B sky130_fd_sc_hd__nand2_1
X_8399_ _8396_/Y _8397_/X _8255_/B _8398_/X VGND VGND VPWR VPWR _8399_/X sky130_fd_sc_hd__a211o_1
X_7419_ _7419_/A _7419_/B _7419_/C _7419_/D VGND VGND VPWR VPWR _7419_/X sky130_fd_sc_hd__and4_1
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput91 _9133_/Q VGND VGND VPWR VPWR F[4] sky130_fd_sc_hd__buf_2
Xoutput80 _9152_/Q VGND VGND VPWR VPWR F[23] sky130_fd_sc_hd__buf_2
XFILLER_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7770_ _7770_/A _8349_/B _7770_/C VGND VGND VPWR VPWR _7771_/B sky130_fd_sc_hd__and3_1
XFILLER_91_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4982_ _4982_/A VGND VGND VPWR VPWR _5743_/S sky130_fd_sc_hd__clkbuf_2
X_6721_ _9209_/Q VGND VGND VPWR VPWR _7307_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6652_ _6652_/A VGND VGND VPWR VPWR _9082_/D sky130_fd_sc_hd__clkbuf_1
X_5603_ _5754_/B _5602_/X _5603_/S VGND VGND VPWR VPWR _5603_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8322_ _8322_/A _8909_/B _8322_/C VGND VGND VPWR VPWR _8423_/B sky130_fd_sc_hd__and3_1
X_6583_ _6719_/A _6719_/B VGND VGND VPWR VPWR _6716_/A sky130_fd_sc_hd__xnor2_2
X_5534_ _5534_/A VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8253_ _8254_/A _8254_/B VGND VGND VPWR VPWR _8255_/A sky130_fd_sc_hd__and2_1
X_5465_ _5141_/A _5179_/A _5464_/X _5219_/X VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__a211o_1
X_8184_ _8054_/A _8184_/B VGND VGND VPWR VPWR _8197_/A sky130_fd_sc_hd__and2b_1
X_7204_ _7204_/A _7204_/B VGND VGND VPWR VPWR _7208_/A sky130_fd_sc_hd__xnor2_1
X_7135_ _7134_/A _7134_/B _7134_/C VGND VGND VPWR VPWR _7235_/A sky130_fd_sc_hd__o21ai_2
X_5396_ _5245_/X _5187_/X _5392_/X _5395_/Y VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7066_ _7066_/A _7066_/B VGND VGND VPWR VPWR _7068_/B sky130_fd_sc_hd__or2_1
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6017_ _6018_/B _6018_/C _6018_/A VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__a21o_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _8093_/A VGND VGND VPWR VPWR _8351_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_42_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7899_ _7782_/A _7899_/B VGND VGND VPWR VPWR _7899_/X sky130_fd_sc_hd__and2b_2
X_6919_ _6919_/A _6803_/B VGND VGND VPWR VPWR _6934_/A sky130_fd_sc_hd__or2b_1
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5250_ _9076_/Q VGND VGND VPWR VPWR _5404_/A sky130_fd_sc_hd__clkinv_2
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5181_ _5181_/A VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8940_ _8902_/A _8902_/B _8890_/B VGND VGND VPWR VPWR _8941_/B sky130_fd_sc_hd__o21ai_1
XFILLER_95_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8871_ _8913_/A _8871_/B VGND VGND VPWR VPWR _8872_/C sky130_fd_sc_hd__or2_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7822_ _7822_/A _7822_/B _7822_/C _7822_/D VGND VGND VPWR VPWR _7944_/A sky130_fd_sc_hd__and4_1
X_7753_ _8069_/A _8091_/D VGND VGND VPWR VPWR _7754_/B sky130_fd_sc_hd__nand2_1
X_4965_ _4550_/A _4962_/X _4963_/Y _4964_/X VGND VGND VPWR VPWR _4965_/X sky130_fd_sc_hd__a2bb2o_1
X_6704_ _6704_/A _6704_/B VGND VGND VPWR VPWR _6706_/A sky130_fd_sc_hd__nor2_1
X_7684_ _7684_/A _7684_/B _7684_/C VGND VGND VPWR VPWR _7686_/B sky130_fd_sc_hd__and3_1
X_4896_ _4896_/A VGND VGND VPWR VPWR _5676_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6635_ _6734_/A _6635_/B VGND VGND VPWR VPWR _6637_/C sky130_fd_sc_hd__or2_2
X_6566_ _6566_/A _6524_/B VGND VGND VPWR VPWR _6580_/B sky130_fd_sc_hd__or2b_1
X_8305_ _8305_/A _8305_/B VGND VGND VPWR VPWR _8307_/B sky130_fd_sc_hd__or2_1
X_5517_ _5215_/X _5634_/A _5515_/X _5516_/Y _5222_/X VGND VGND VPWR VPWR _5517_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8236_ _8161_/B _8236_/B VGND VGND VPWR VPWR _8236_/X sky130_fd_sc_hd__and2b_1
X_6497_ _7730_/B VGND VGND VPWR VPWR _7962_/B sky130_fd_sc_hd__buf_2
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5448_ _5245_/A _5403_/X _5446_/X _5447_/Y _5391_/X VGND VGND VPWR VPWR _5448_/X
+ sky130_fd_sc_hd__a221o_1
X_8167_ _8166_/A _8166_/B _8166_/C VGND VGND VPWR VPWR _8168_/C sky130_fd_sc_hd__o21ai_4
X_5379_ _4600_/A _5212_/X _5378_/X VGND VGND VPWR VPWR _5379_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8098_ _8098_/A _8098_/B VGND VGND VPWR VPWR _8166_/B sky130_fd_sc_hd__and2_1
X_7118_ _7118_/A _7988_/B VGND VGND VPWR VPWR _7122_/A sky130_fd_sc_hd__nand2_1
X_7049_ _7048_/A _7048_/B _7048_/C VGND VGND VPWR VPWR _7104_/A sky130_fd_sc_hd__a21o_2
XFILLER_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4750_ _4816_/A _4750_/B VGND VGND VPWR VPWR _4842_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ _9122_/Q _9114_/Q VGND VGND VPWR VPWR _4691_/B sky130_fd_sc_hd__xor2_1
X_6420_ _6341_/A _6340_/A _6340_/B VGND VGND VPWR VPWR _6489_/A sky130_fd_sc_hd__o21ba_2
X_6351_ _6260_/A _6351_/B VGND VGND VPWR VPWR _6367_/A sky130_fd_sc_hd__and2b_1
X_5302_ _5403_/A _5122_/X _5300_/X _5301_/Y VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__a22o_1
X_9070_ _9090_/CLK _9070_/D VGND VGND VPWR VPWR _9070_/Q sky130_fd_sc_hd__dfxtp_2
X_6282_ _6282_/A _6282_/B VGND VGND VPWR VPWR _6283_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8021_ _8128_/A VGND VGND VPWR VPWR _8024_/A sky130_fd_sc_hd__inv_2
X_5233_ _5736_/S VGND VGND VPWR VPWR _5572_/S sky130_fd_sc_hd__buf_2
X_5164_ _5164_/A VGND VGND VPWR VPWR _5367_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _5093_/Y _4998_/A _5041_/A _5741_/S VGND VGND VPWR VPWR _5095_/X sky130_fd_sc_hd__a31o_1
X_8923_ _8923_/A VGND VGND VPWR VPWR _8957_/A sky130_fd_sc_hd__inv_2
XFILLER_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8854_ _8855_/A _8855_/B VGND VGND VPWR VPWR _8856_/A sky130_fd_sc_hd__nand2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7805_ _7805_/A _7805_/B VGND VGND VPWR VPWR _7902_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8785_ _8785_/A _8836_/B VGND VGND VPWR VPWR _8787_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5997_ _5997_/A _5997_/B _5997_/C VGND VGND VPWR VPWR _5999_/A sky130_fd_sc_hd__nand3_1
X_7736_ _7736_/A _7736_/B VGND VGND VPWR VPWR _7843_/B sky130_fd_sc_hd__xnor2_1
X_4948_ _4845_/Y _4920_/A _4947_/Y VGND VGND VPWR VPWR _4948_/Y sky130_fd_sc_hd__a21oi_1
X_7667_ _7683_/A _7667_/B VGND VGND VPWR VPWR _7668_/C sky130_fd_sc_hd__xnor2_1
XFILLER_20_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4879_ _5177_/A VGND VGND VPWR VPWR _4880_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6618_ _6716_/A _6716_/B _6716_/C VGND VGND VPWR VPWR _6618_/X sky130_fd_sc_hd__or3_1
X_7598_ _7684_/B _7684_/C VGND VGND VPWR VPWR _7599_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_6549_ _6548_/B _6548_/C _6548_/A VGND VGND VPWR VPWR _6550_/B sky130_fd_sc_hd__o21a_1
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8219_ _8219_/A _8219_/B VGND VGND VPWR VPWR _8221_/A sky130_fd_sc_hd__nor2_1
X_9199_ _9199_/CLK _9199_/D VGND VGND VPWR VPWR _9199_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5920_ _7361_/C VGND VGND VPWR VPWR _7767_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5851_ _6169_/A _9194_/Q VGND VGND VPWR VPWR _5854_/B sky130_fd_sc_hd__nand2_1
X_8570_ _8571_/A _8571_/B _8571_/C VGND VGND VPWR VPWR _8570_/Y sky130_fd_sc_hd__o21ai_2
X_5782_ _4541_/X _5781_/X _5741_/S VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__o21a_1
X_4802_ _4770_/X _4764_/X _4801_/X _5187_/A VGND VGND VPWR VPWR _4802_/X sky130_fd_sc_hd__a211o_1
X_7521_ _7521_/A _7661_/A VGND VGND VPWR VPWR _7522_/C sky130_fd_sc_hd__nor2_1
X_4733_ _9107_/Q VGND VGND VPWR VPWR _5738_/S sky130_fd_sc_hd__inv_2
X_7452_ _7452_/A _7355_/B VGND VGND VPWR VPWR _7474_/B sky130_fd_sc_hd__or2b_1
X_6403_ _7152_/A VGND VGND VPWR VPWR _6927_/C sky130_fd_sc_hd__clkbuf_2
X_4664_ _5222_/A VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__clkbuf_2
X_7383_ _7383_/A _7383_/B VGND VGND VPWR VPWR _7384_/B sky130_fd_sc_hd__nand2_2
X_4595_ _9099_/Q VGND VGND VPWR VPWR _5002_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9122_ _9222_/CLK hold7/X VGND VGND VPWR VPWR _9122_/Q sky130_fd_sc_hd__dfxtp_2
X_6334_ _6259_/A _6258_/A _6258_/B VGND VGND VPWR VPWR _6345_/A sky130_fd_sc_hd__o21ba_2
X_9053_ _9052_/A _9052_/C _6053_/B _9052_/Y VGND VGND VPWR VPWR _9074_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6265_ _6262_/Y _6263_/X _6264_/C _6264_/Y VGND VGND VPWR VPWR _6288_/B sky130_fd_sc_hd__o211ai_2
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8004_ _7894_/A _7894_/B _7893_/B VGND VGND VPWR VPWR _8005_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5216_ _5144_/A _5150_/Y _4846_/A VGND VGND VPWR VPWR _5216_/Y sky130_fd_sc_hd__a21oi_1
X_6196_ _6361_/C VGND VGND VPWR VPWR _8091_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5147_ _9068_/Q _5146_/X _4847_/X VGND VGND VPWR VPWR _5147_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5078_ _5070_/X _5075_/X _5076_/X _5077_/Y _4726_/X VGND VGND VPWR VPWR _5078_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8906_ _8906_/A _8849_/A VGND VGND VPWR VPWR _8907_/A sky130_fd_sc_hd__or2b_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8837_ _8889_/A _8837_/B VGND VGND VPWR VPWR _8839_/B sky130_fd_sc_hd__and2_1
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8768_ _8768_/A _8768_/B _8766_/Y VGND VGND VPWR VPWR _8768_/X sky130_fd_sc_hd__or3b_1
XFILLER_25_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7719_ _7717_/X _7718_/Y _7621_/C _7622_/B VGND VGND VPWR VPWR _7724_/B sky130_fd_sc_hd__o211ai_1
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8699_ _8699_/A _8699_/B VGND VGND VPWR VPWR _8701_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6048_/A _6049_/C _9052_/C _9052_/A VGND VGND VPWR VPWR _6051_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5001_ _5001_/A VGND VGND VPWR VPWR _5164_/A sky130_fd_sc_hd__clkbuf_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6952_ _6952_/A _6952_/B VGND VGND VPWR VPWR _6952_/X sky130_fd_sc_hd__or2_1
X_6883_ _6883_/A _6793_/A VGND VGND VPWR VPWR _6901_/A sky130_fd_sc_hd__or2b_1
X_5903_ _5903_/A _5903_/B _5903_/C VGND VGND VPWR VPWR _5906_/B sky130_fd_sc_hd__nand3_1
X_8622_ _8622_/A _8622_/B VGND VGND VPWR VPWR _8624_/C sky130_fd_sc_hd__or2_1
X_5834_ _5834_/A _5834_/B VGND VGND VPWR VPWR _5883_/B sky130_fd_sc_hd__xor2_1
X_8553_ _8554_/A _8554_/B VGND VGND VPWR VPWR _8556_/B sky130_fd_sc_hd__nand2_1
X_5765_ _5765_/A _5765_/B _5765_/C VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__or3_1
X_7504_ _7643_/A _7501_/Y _7635_/A VGND VGND VPWR VPWR _7513_/A sky130_fd_sc_hd__a21o_1
X_8484_ _8481_/Y _8482_/X _8479_/Y _8480_/X VGND VGND VPWR VPWR _8565_/A sky130_fd_sc_hd__o211a_2
X_5696_ _5606_/A _5695_/X _5696_/S VGND VGND VPWR VPWR _5696_/X sky130_fd_sc_hd__mux2_1
X_4716_ _4716_/A VGND VGND VPWR VPWR _4717_/S sky130_fd_sc_hd__clkbuf_2
X_7435_ _7435_/A _7583_/A _7706_/C _7583_/D VGND VGND VPWR VPWR _7436_/B sky130_fd_sc_hd__and4_1
X_4647_ _4846_/A VGND VGND VPWR VPWR _4856_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7366_ _7259_/A _7259_/D _9182_/Q _7119_/B VGND VGND VPWR VPWR _7368_/A sky130_fd_sc_hd__a22oi_2
X_6317_ _6663_/C VGND VGND VPWR VPWR _7938_/B sky130_fd_sc_hd__clkbuf_2
X_9105_ _9116_/CLK _9105_/D VGND VGND VPWR VPWR _9105_/Q sky130_fd_sc_hd__dfxtp_2
X_4578_ _5252_/A _5286_/A VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7297_ _7189_/C _7696_/B _7189_/D _7187_/X VGND VGND VPWR VPWR _7298_/B sky130_fd_sc_hd__a31o_1
X_9036_ _9035_/A _9035_/B _9035_/C VGND VGND VPWR VPWR _9036_/X sky130_fd_sc_hd__a21o_1
X_6248_ _6248_/A _6332_/B _6248_/C VGND VGND VPWR VPWR _6263_/C sky130_fd_sc_hd__nand3_1
XFILLER_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6179_ _6179_/A _6179_/B VGND VGND VPWR VPWR _6180_/B sky130_fd_sc_hd__xnor2_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5550_ _4566_/X _5020_/X _4697_/A VGND VGND VPWR VPWR _5550_/Y sky130_fd_sc_hd__a21oi_1
X_5481_ _5433_/X _5480_/X _5481_/S VGND VGND VPWR VPWR _5481_/X sky130_fd_sc_hd__mux2_1
XANTENNA_0 _9180_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7220_ _7694_/B _7730_/B VGND VGND VPWR VPWR _7224_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7151_ _7152_/B _7042_/D _7330_/A _7042_/B VGND VGND VPWR VPWR _7151_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7082_ _6500_/B _6825_/C _7706_/D _6405_/B VGND VGND VPWR VPWR _7084_/A sky130_fd_sc_hd__a22oi_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6187_/A _6102_/B VGND VGND VPWR VPWR _6104_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6107_/A _6107_/B VGND VGND VPWR VPWR _6108_/B sky130_fd_sc_hd__xor2_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7984_ _7984_/A _7997_/A VGND VGND VPWR VPWR _7993_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6935_ _6934_/A _6934_/B _6934_/C VGND VGND VPWR VPWR _6988_/A sky130_fd_sc_hd__a21o_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6866_ _6830_/A _6830_/B _6865_/X VGND VGND VPWR VPWR _6868_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8605_ _8518_/A _8520_/B _8518_/B VGND VGND VPWR VPWR _8661_/A sky130_fd_sc_hd__o21ba_1
X_6797_ _6665_/A _6664_/A _6664_/B VGND VGND VPWR VPWR _6919_/A sky130_fd_sc_hd__o21ba_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5817_ _9195_/Q VGND VGND VPWR VPWR _6055_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8536_ _8639_/A _8898_/B VGND VGND VPWR VPWR _8537_/B sky130_fd_sc_hd__nand2_1
X_5748_ _5339_/A _5746_/X _5747_/Y _5450_/X _5618_/X VGND VGND VPWR VPWR _5749_/B
+ sky130_fd_sc_hd__o221a_1
X_8467_ _8467_/A VGND VGND VPWR VPWR _8666_/A sky130_fd_sc_hd__clkbuf_2
X_5679_ _4940_/A _5389_/A _9094_/Q VGND VGND VPWR VPWR _5679_/Y sky130_fd_sc_hd__a21oi_1
X_8398_ _8256_/A _8398_/B VGND VGND VPWR VPWR _8398_/X sky130_fd_sc_hd__and2b_1
X_7418_ _7421_/D VGND VGND VPWR VPWR _7418_/Y sky130_fd_sc_hd__clkinv_2
X_7349_ _7349_/A _9200_/Q _9177_/Q _9178_/Q VGND VGND VPWR VPWR _7349_/X sky130_fd_sc_hd__and4_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9019_ _9038_/A _9038_/B VGND VGND VPWR VPWR _9022_/A sky130_fd_sc_hd__xnor2_2
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput70 _9143_/Q VGND VGND VPWR VPWR F[14] sky130_fd_sc_hd__buf_2
Xoutput92 _9134_/Q VGND VGND VPWR VPWR F[5] sky130_fd_sc_hd__buf_2
XFILLER_95_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput81 _9153_/Q VGND VGND VPWR VPWR F[24] sky130_fd_sc_hd__buf_2
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _4980_/A _4978_/Y _4979_/X _4980_/Y _4930_/A VGND VGND VPWR VPWR _4981_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6720_ _7299_/A _8519_/A _6571_/A _6569_/A VGND VGND VPWR VPWR _6730_/A sky130_fd_sc_hd__a31o_1
XFILLER_44_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6651_ _6651_/A _6654_/B VGND VGND VPWR VPWR _6652_/A sky130_fd_sc_hd__and2_1
X_5602_ _5534_/X _5601_/X _5674_/S VGND VGND VPWR VPWR _5602_/X sky130_fd_sc_hd__mux2_1
X_6582_ _6582_/A _6737_/A VGND VGND VPWR VPWR _6719_/B sky130_fd_sc_hd__nand2_1
X_8321_ _8322_/A _8816_/B _8322_/C VGND VGND VPWR VPWR _8323_/A sky130_fd_sc_hd__a21oi_1
X_5533_ _5509_/X _5510_/X _5511_/X _5531_/X _5532_/X VGND VGND VPWR VPWR _9140_/D
+ sky130_fd_sc_hd__o221a_4
XFILLER_105_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8252_ _8252_/A _8252_/B VGND VGND VPWR VPWR _8254_/B sky130_fd_sc_hd__xnor2_1
X_5464_ _4570_/A _5246_/Y _5462_/Y _5463_/X _5251_/A VGND VGND VPWR VPWR _5464_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8183_ _8183_/A _8183_/B VGND VGND VPWR VPWR _8201_/A sky130_fd_sc_hd__xor2_1
X_7203_ _7203_/A _7313_/B VGND VGND VPWR VPWR _7204_/B sky130_fd_sc_hd__xnor2_1
X_5395_ _5394_/X _5276_/X _5105_/A VGND VGND VPWR VPWR _5395_/Y sky130_fd_sc_hd__a21oi_1
X_7134_ _7134_/A _7134_/B _7134_/C VGND VGND VPWR VPWR _7136_/A sky130_fd_sc_hd__or3_1
XFILLER_86_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7065_ _7065_/A _7066_/B VGND VGND VPWR VPWR _9086_/D sky130_fd_sc_hd__xnor2_1
X_6016_ _6016_/A _6016_/B VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _7967_/A _7967_/B VGND VGND VPWR VPWR _7970_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7898_ _7898_/A _7898_/B VGND VGND VPWR VPWR _7901_/A sky130_fd_sc_hd__xor2_2
XFILLER_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6918_ _6766_/A _6766_/B _6917_/X VGND VGND VPWR VPWR _6961_/A sky130_fd_sc_hd__a21oi_1
X_6849_ _6849_/A _6952_/B VGND VGND VPWR VPWR _9084_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8519_ _8519_/A _8664_/C VGND VGND VPWR VPWR _8520_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5180_ _5177_/X _5179_/X _5126_/A VGND VGND VPWR VPWR _5180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8870_ _8870_/A _8870_/B VGND VGND VPWR VPWR _8871_/B sky130_fd_sc_hd__and2_1
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7821_ _7938_/A _7706_/C _7583_/D _7706_/B VGND VGND VPWR VPWR _7823_/A sky130_fd_sc_hd__a22oi_1
XFILLER_64_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7752_ _8071_/A _8156_/C VGND VGND VPWR VPWR _7752_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4964_ _4963_/A _4963_/B _5129_/A VGND VGND VPWR VPWR _4964_/X sky130_fd_sc_hd__o21a_1
X_6703_ _7307_/B _7042_/B _6572_/D _7307_/A VGND VGND VPWR VPWR _6704_/B sky130_fd_sc_hd__a22oi_2
X_7683_ _7683_/A _7667_/B VGND VGND VPWR VPWR _7788_/B sky130_fd_sc_hd__or2b_1
X_4895_ _5336_/S _4893_/Y _4894_/X VGND VGND VPWR VPWR _4895_/X sky130_fd_sc_hd__a21o_1
X_6634_ _6632_/C _6831_/A VGND VGND VPWR VPWR _6635_/B sky130_fd_sc_hd__and2b_1
X_6565_ _6565_/A _6565_/B _6611_/B VGND VGND VPWR VPWR _6580_/A sky130_fd_sc_hd__or3_1
X_8304_ _8304_/A _8304_/B VGND VGND VPWR VPWR _8305_/B sky130_fd_sc_hd__nor2_1
X_5516_ _4862_/A _9084_/Q _5215_/A VGND VGND VPWR VPWR _5516_/Y sky130_fd_sc_hd__a21oi_1
X_6496_ _9207_/Q VGND VGND VPWR VPWR _7730_/B sky130_fd_sc_hd__clkbuf_2
X_8235_ _8220_/A _9004_/B _8221_/A _8219_/B VGND VGND VPWR VPWR _8336_/A sky130_fd_sc_hd__a31oi_2
X_5447_ _5394_/X _5126_/X _5181_/X VGND VGND VPWR VPWR _5447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8166_ _8166_/A _8166_/B _8166_/C VGND VGND VPWR VPWR _8168_/B sky130_fd_sc_hd__or3_1
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5378_ _5378_/A VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__clkbuf_2
X_8097_ _8098_/A _8098_/B VGND VGND VPWR VPWR _8099_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7117_ _7117_/A _7246_/B VGND VGND VPWR VPWR _7251_/A sky130_fd_sc_hd__nor2_1
X_7048_ _7048_/A _7048_/B _7048_/C VGND VGND VPWR VPWR _7050_/A sky130_fd_sc_hd__nand3_1
XFILLER_47_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8999_ _8999_/A _8999_/B VGND VGND VPWR VPWR _9001_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4680_ _4691_/A _4680_/B VGND VGND VPWR VPWR _9152_/D sky130_fd_sc_hd__xnor2_4
X_6350_ _6350_/A _6350_/B _6350_/C VGND VGND VPWR VPWR _6372_/C sky130_fd_sc_hd__and3_1
X_5301_ _5271_/A _5189_/X _5181_/A VGND VGND VPWR VPWR _5301_/Y sky130_fd_sc_hd__a21oi_1
X_6281_ _6282_/A _6282_/B VGND VGND VPWR VPWR _6370_/A sky130_fd_sc_hd__and2_1
XFILLER_102_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8020_ _8020_/A _8020_/B VGND VGND VPWR VPWR _8128_/A sky130_fd_sc_hd__nor2_1
X_5232_ _4726_/X _5212_/X _5231_/X VGND VGND VPWR VPWR _5232_/Y sky130_fd_sc_hd__o21ai_1
X_5163_ _5136_/X _5482_/A _5159_/X _5162_/Y _4558_/A VGND VGND VPWR VPWR _5163_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5094_ _5093_/Y _5028_/A _5041_/A VGND VGND VPWR VPWR _5094_/Y sky130_fd_sc_hd__a21oi_1
X_8922_ _8965_/A _8922_/B VGND VGND VPWR VPWR _9106_/D sky130_fd_sc_hd__xnor2_1
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8853_ _8853_/A _8907_/B VGND VGND VPWR VPWR _8855_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7804_ _7804_/A _7804_/B VGND VGND VPWR VPWR _7805_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8784_ _8784_/A _8784_/B VGND VGND VPWR VPWR _8836_/B sky130_fd_sc_hd__and2_1
XFILLER_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5996_ _5993_/X _5994_/Y _5930_/B _5930_/Y VGND VGND VPWR VPWR _5997_/C sky130_fd_sc_hd__o211ai_1
X_7735_ _8093_/A _8290_/A VGND VGND VPWR VPWR _7736_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4947_ _4845_/Y _4920_/A _5215_/A VGND VGND VPWR VPWR _4947_/Y sky130_fd_sc_hd__o21ai_1
X_7666_ _7666_/A _7682_/A VGND VGND VPWR VPWR _7667_/B sky130_fd_sc_hd__xnor2_1
X_4878_ _4878_/A VGND VGND VPWR VPWR _5177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6617_ _6616_/A _6616_/B _6616_/C VGND VGND VPWR VPWR _6716_/C sky130_fd_sc_hd__a21oi_4
X_7597_ _7686_/A VGND VGND VPWR VPWR _7684_/C sky130_fd_sc_hd__inv_2
XFILLER_20_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6548_ _6548_/A _6548_/B _6548_/C VGND VGND VPWR VPWR _6550_/A sky130_fd_sc_hd__nor3_1
X_6479_ _6479_/A VGND VGND VPWR VPWR _9080_/D sky130_fd_sc_hd__clkbuf_1
X_8218_ _8217_/A _8217_/B _8216_/Y VGND VGND VPWR VPWR _8219_/B sky130_fd_sc_hd__o21ba_1
X_9198_ _9216_/CLK _9198_/D VGND VGND VPWR VPWR _9198_/Q sky130_fd_sc_hd__dfxtp_2
X_8149_ _8337_/A _8464_/B _8542_/C _8517_/A VGND VGND VPWR VPWR _8151_/A sky130_fd_sc_hd__a22oi_1
XFILLER_59_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5850_ _9166_/Q VGND VGND VPWR VPWR _6169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5781_ _5632_/A _5780_/X _5305_/S VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__o21a_1
X_4801_ _5403_/A _4798_/X _4799_/Y _5671_/S VGND VGND VPWR VPWR _4801_/X sky130_fd_sc_hd__o211a_1
X_7520_ _7518_/C _7518_/Y _7658_/B _7517_/X VGND VGND VPWR VPWR _7661_/A sky130_fd_sc_hd__a211oi_4
X_4732_ _4698_/X _4731_/X _5354_/S VGND VGND VPWR VPWR _4732_/X sky130_fd_sc_hd__mux2_1
X_7451_ _7317_/B _7449_/X _7447_/X _7559_/A VGND VGND VPWR VPWR _7559_/B sky130_fd_sc_hd__a211oi_2
X_4663_ _4789_/A VGND VGND VPWR VPWR _5222_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6402_ _7295_/C _7462_/A VGND VGND VPWR VPWR _6407_/A sky130_fd_sc_hd__nand2_1
X_7382_ _7382_/A _7382_/B VGND VGND VPWR VPWR _7528_/A sky130_fd_sc_hd__nand2_2
X_4594_ _4566_/X _4588_/X _5432_/A VGND VGND VPWR VPWR _4594_/X sky130_fd_sc_hd__a21o_1
X_9121_ _9223_/CLK hold16/X VGND VGND VPWR VPWR _9121_/Q sky130_fd_sc_hd__dfxtp_2
X_6333_ _6332_/A _6332_/B _6332_/C VGND VGND VPWR VPWR _6347_/C sky130_fd_sc_hd__a21o_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9052_ _9052_/A _9052_/B _9052_/C VGND VGND VPWR VPWR _9052_/Y sky130_fd_sc_hd__nand3_1
X_6264_ _6264_/A _6264_/B _6264_/C VGND VGND VPWR VPWR _6264_/Y sky130_fd_sc_hd__nand3_1
X_8003_ _8003_/A _8003_/B VGND VGND VPWR VPWR _8005_/A sky130_fd_sc_hd__xor2_2
X_5215_ _5215_/A VGND VGND VPWR VPWR _5215_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X VGND VGND VPWR VPWR _9210_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6195_ _6828_/A VGND VGND VPWR VPWR _6968_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5146_ _5146_/A VGND VGND VPWR VPWR _5146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5077_ _4963_/A _5046_/Y _5173_/A VGND VGND VPWR VPWR _5077_/Y sky130_fd_sc_hd__o21ai_1
X_8905_ _8947_/A _8905_/B VGND VGND VPWR VPWR _8923_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8836_ _8836_/A _8836_/B _8836_/C VGND VGND VPWR VPWR _8837_/B sky130_fd_sc_hd__or3_1
XFILLER_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8767_ _8768_/A _8768_/B _8766_/Y VGND VGND VPWR VPWR _8769_/A sky130_fd_sc_hd__o21ba_1
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5979_ _5979_/A _5979_/B _5979_/C VGND VGND VPWR VPWR _6037_/A sky130_fd_sc_hd__nand3_2
X_7718_ _7718_/A _7718_/B VGND VGND VPWR VPWR _7718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8698_ _8624_/X _8627_/A _8697_/C VGND VGND VPWR VPWR _8699_/B sky130_fd_sc_hd__o21ba_1
X_7649_ _7770_/A _8243_/B _9184_/Q _7647_/A VGND VGND VPWR VPWR _7649_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A VGND VGND VPWR VPWR clkbuf_4_9_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_6951_ _6957_/A _6957_/B VGND VGND VPWR VPWR _7066_/A sky130_fd_sc_hd__xnor2_1
X_6882_ _6882_/A _6882_/B _6882_/C _6960_/A VGND VGND VPWR VPWR _6960_/B sky130_fd_sc_hd__nor4_1
X_5902_ _5903_/B _5903_/C _5903_/A VGND VGND VPWR VPWR _5906_/A sky130_fd_sc_hd__a21o_1
X_8621_ _8622_/A _8622_/B VGND VGND VPWR VPWR _8624_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ _5833_/A _5898_/C VGND VGND VPWR VPWR _5883_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8552_ _8552_/A _8552_/B VGND VGND VPWR VPWR _8554_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7503_ _7767_/A _8091_/D _7503_/C VGND VGND VPWR VPWR _7635_/A sky130_fd_sc_hd__and3_1
X_5764_ _5281_/S _5763_/X _4687_/X _4541_/X VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__a211o_1
X_8483_ _8479_/Y _8480_/X _8481_/Y _8482_/X VGND VGND VPWR VPWR _8483_/Y sky130_fd_sc_hd__a211oi_2
X_4715_ _5000_/A VGND VGND VPWR VPWR _4716_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5695_ _5754_/A _5694_/X _5695_/S VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__mux2_1
X_7434_ _6679_/A _7938_/C _8050_/D _7694_/B VGND VGND VPWR VPWR _7436_/A sky130_fd_sc_hd__a22oi_1
X_4646_ _4783_/A VGND VGND VPWR VPWR _4846_/A sky130_fd_sc_hd__clkbuf_2
X_7365_ _7365_/A _7986_/B VGND VGND VPWR VPWR _7369_/A sky130_fd_sc_hd__nand2_1
X_4577_ _4776_/A VGND VGND VPWR VPWR _5286_/A sky130_fd_sc_hd__clkbuf_2
X_6316_ _9174_/Q VGND VGND VPWR VPWR _6663_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_9104_ _9116_/CLK _9104_/D VGND VGND VPWR VPWR _9104_/Q sky130_fd_sc_hd__dfxtp_2
X_7296_ _7296_/A _7296_/B VGND VGND VPWR VPWR _7298_/A sky130_fd_sc_hd__nor2_1
X_9035_ _9035_/A _9035_/B _9035_/C VGND VGND VPWR VPWR _9037_/A sky130_fd_sc_hd__and3_1
X_6247_ _6248_/A _6332_/B _6248_/C VGND VGND VPWR VPWR _6263_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6178_ _6567_/B _6607_/B VGND VGND VPWR VPWR _6179_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5129_ _5129_/A VGND VGND VPWR VPWR _5129_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8819_ _8819_/A _8819_/B _8819_/C VGND VGND VPWR VPWR _8821_/A sky130_fd_sc_hd__nor3_1
XFILLER_13_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5480_ _5402_/X _5479_/X _5553_/S VGND VGND VPWR VPWR _5480_/X sky130_fd_sc_hd__mux2_1
XANTENNA_1 _9180_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7150_ _7150_/A _7150_/B VGND VGND VPWR VPWR _7159_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7081_ _7081_/A _9210_/Q VGND VGND VPWR VPWR _7085_/A sky130_fd_sc_hd__nand2_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6186_/A _6101_/B VGND VGND VPWR VPWR _6102_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6032_/A _6032_/B VGND VGND VPWR VPWR _6107_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7983_ _8137_/A _8717_/A _7874_/A _7870_/X VGND VGND VPWR VPWR _7995_/A sky130_fd_sc_hd__a31o_1
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6934_ _6934_/A _6934_/B _6934_/C VGND VGND VPWR VPWR _6936_/A sky130_fd_sc_hd__nand3_1
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8604_ _8604_/A _8604_/B VGND VGND VPWR VPWR _8622_/A sky130_fd_sc_hd__or2_1
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _6830_/A _6830_/B _6832_/A VGND VGND VPWR VPWR _6865_/X sky130_fd_sc_hd__o21a_1
X_6796_ _6795_/A _6795_/B _6795_/C VGND VGND VPWR VPWR _6808_/C sky130_fd_sc_hd__a21o_1
X_5816_ _6859_/B VGND VGND VPWR VPWR _6361_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8535_ _8633_/B _8535_/B VGND VGND VPWR VPWR _8537_/A sky130_fd_sc_hd__xnor2_2
XFILLER_10_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5747_ _5200_/A _5558_/X _4650_/A VGND VGND VPWR VPWR _5747_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8466_ _8466_/A VGND VGND VPWR VPWR _8538_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7417_ _7199_/A _9211_/Q _9212_/Q _7083_/A VGND VGND VPWR VPWR _7421_/D sky130_fd_sc_hd__a22o_1
X_5678_ _5678_/A VGND VGND VPWR VPWR _5765_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_8397_ _8397_/A _8397_/B VGND VGND VPWR VPWR _8397_/X sky130_fd_sc_hd__or2_2
X_4629_ _4629_/A _9109_/Q _9110_/Q _9112_/Q VGND VGND VPWR VPWR _4677_/A sky130_fd_sc_hd__or4_1
XFILLER_104_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7348_ _7348_/A _7348_/B VGND VGND VPWR VPWR _7490_/A sky130_fd_sc_hd__nand2_1
X_7279_ _7168_/Y _7171_/B _7276_/X _7277_/Y VGND VGND VPWR VPWR _7284_/C sky130_fd_sc_hd__a211o_1
X_9018_ _9018_/A _8996_/X VGND VGND VPWR VPWR _9038_/B sky130_fd_sc_hd__or2b_1
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput82 _9154_/Q VGND VGND VPWR VPWR F[25] sky130_fd_sc_hd__buf_2
Xoutput93 _9135_/Q VGND VGND VPWR VPWR F[6] sky130_fd_sc_hd__buf_2
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput71 _9144_/Q VGND VGND VPWR VPWR F[15] sky130_fd_sc_hd__buf_2
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4980_ _4980_/A _4980_/B VGND VGND VPWR VPWR _4980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6650_ _6649_/A _6649_/B _6649_/C VGND VGND VPWR VPWR _6654_/B sky130_fd_sc_hd__o21ai_1
X_5601_ _5509_/X _5600_/X _5673_/S VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__mux2_1
X_6581_ _6580_/A _6580_/B _6580_/C VGND VGND VPWR VPWR _6737_/A sky130_fd_sc_hd__a21o_1
X_8320_ _8320_/A _8423_/A VGND VGND VPWR VPWR _8322_/C sky130_fd_sc_hd__nor2_1
X_5532_ _5532_/A _5604_/B VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__or2_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8251_ _8251_/A _8361_/A VGND VGND VPWR VPWR _8252_/B sky130_fd_sc_hd__xnor2_1
X_5463_ _4849_/A _5172_/A _5146_/A _5166_/Y _4783_/X VGND VGND VPWR VPWR _5463_/X
+ sky130_fd_sc_hd__a221o_1
X_8182_ _8322_/A _8798_/B VGND VGND VPWR VPWR _8183_/B sky130_fd_sc_hd__nand2_1
X_7202_ _7202_/A _7202_/B VGND VGND VPWR VPWR _7313_/B sky130_fd_sc_hd__xnor2_1
X_5394_ _5394_/A VGND VGND VPWR VPWR _5394_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7133_ _7133_/A _7133_/B VGND VGND VPWR VPWR _7134_/C sky130_fd_sc_hd__xnor2_1
XFILLER_86_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7064_ _7064_/A _7064_/B VGND VGND VPWR VPWR _7066_/B sky130_fd_sc_hd__xor2_1
XFILLER_100_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6015_ _6859_/A _7254_/C VGND VGND VPWR VPWR _6016_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _8156_/A _8156_/B _8148_/A _7966_/D VGND VGND VPWR VPWR _7967_/B sky130_fd_sc_hd__and4_1
X_7897_ _7897_/A _8009_/B VGND VGND VPWR VPWR _7898_/B sky130_fd_sc_hd__xnor2_4
X_6917_ _6765_/B _6917_/B VGND VGND VPWR VPWR _6917_/X sky130_fd_sc_hd__and2b_1
XFILLER_35_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6848_ _6848_/A _6848_/B VGND VGND VPWR VPWR _6952_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8518_ _8518_/A _8518_/B VGND VGND VPWR VPWR _8520_/A sky130_fd_sc_hd__nor2_1
X_6779_ _6590_/B _7465_/A _7360_/A _7016_/A VGND VGND VPWR VPWR _6780_/B sky130_fd_sc_hd__a22oi_1
X_8449_ _8597_/A _8450_/C _8450_/D _8527_/A VGND VGND VPWR VPWR _8451_/A sky130_fd_sc_hd__a22oi_1
XFILLER_89_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7820_ _7729_/A _7731_/B _7729_/B VGND VGND VPWR VPWR _7826_/A sky130_fd_sc_hd__o21ba_1
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7751_ _7747_/X _8677_/A _7633_/A _7629_/Y VGND VGND VPWR VPWR _7763_/A sky130_fd_sc_hd__a31o_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4963_ _4963_/A _4963_/B VGND VGND VPWR VPWR _4963_/Y sky130_fd_sc_hd__nand2_1
X_6702_ _6702_/A _6702_/B _7152_/A _7042_/D VGND VGND VPWR VPWR _6704_/A sky130_fd_sc_hd__and4_1
X_7682_ _7682_/A _7666_/A VGND VGND VPWR VPWR _7788_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4894_ _4535_/X _4838_/Y _4896_/A VGND VGND VPWR VPWR _4894_/X sky130_fd_sc_hd__a21o_1
X_6633_ _6968_/B _8190_/C VGND VGND VPWR VPWR _6831_/A sky130_fd_sc_hd__nand2_1
X_6564_ _6507_/A _6507_/B _6563_/X VGND VGND VPWR VPWR _6719_/A sky130_fd_sc_hd__a21oi_2
X_8303_ _8304_/A _8304_/B VGND VGND VPWR VPWR _8305_/A sky130_fd_sc_hd__and2_1
X_5515_ _5141_/A _5184_/A _5514_/Y _5219_/X VGND VGND VPWR VPWR _5515_/X sky130_fd_sc_hd__a211o_1
X_6495_ _6493_/X _6495_/B VGND VGND VPWR VPWR _6499_/A sky130_fd_sc_hd__and2b_1
XFILLER_105_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8234_ _8234_/A _8234_/B VGND VGND VPWR VPWR _8331_/B sky130_fd_sc_hd__and2_1
X_5446_ _5177_/X _5117_/A _5444_/X _5445_/Y _4545_/A VGND VGND VPWR VPWR _5446_/X
+ sky130_fd_sc_hd__a221o_1
X_8165_ _8165_/A _8165_/B VGND VGND VPWR VPWR _8166_/C sky130_fd_sc_hd__and2_1
X_5377_ _4667_/A _5604_/A _5375_/X _5376_/Y _5136_/X VGND VGND VPWR VPWR _5377_/X
+ sky130_fd_sc_hd__a221o_1
X_8096_ _8146_/B _8096_/B VGND VGND VPWR VPWR _8098_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7116_ _7246_/A _7114_/Y _7254_/C _7116_/D VGND VGND VPWR VPWR _7246_/B sky130_fd_sc_hd__and4bb_1
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7047_ _7047_/A _7047_/B VGND VGND VPWR VPWR _7048_/C sky130_fd_sc_hd__xnor2_1
XFILLER_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8998_ _8995_/Y _8996_/X _8958_/B _8973_/X VGND VGND VPWR VPWR _8999_/B sky130_fd_sc_hd__a211oi_2
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _7950_/A _7950_/B VGND VGND VPWR VPWR _7951_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5300_ _5177_/A _5124_/X _5298_/X _5299_/Y _5125_/A VGND VGND VPWR VPWR _5300_/X
+ sky130_fd_sc_hd__a221o_1
X_6280_ _6280_/A _6280_/B VGND VGND VPWR VPWR _6282_/B sky130_fd_sc_hd__xnor2_1
X_5231_ _4721_/X _5179_/X _5228_/X _5229_/Y _5230_/X VGND VGND VPWR VPWR _5231_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5162_ _5160_/X _5370_/A _4599_/A VGND VGND VPWR VPWR _5162_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5093_ _5093_/A VGND VGND VPWR VPWR _5093_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8921_ _8921_/A _8921_/B VGND VGND VPWR VPWR _8922_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8852_ _8852_/A _8852_/B VGND VGND VPWR VPWR _8907_/B sky130_fd_sc_hd__nand2_1
X_8783_ _8784_/A _8784_/B VGND VGND VPWR VPWR _8785_/A sky130_fd_sc_hd__nor2_1
X_7803_ _7803_/A _7803_/B VGND VGND VPWR VPWR _7805_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7734_ _7734_/A _7734_/B VGND VGND VPWR VPWR _7736_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5995_ _5930_/B _5930_/Y _5993_/X _5994_/Y VGND VGND VPWR VPWR _5997_/B sky130_fd_sc_hd__a211o_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4946_ _5219_/A _4916_/X _4931_/X _4945_/X VGND VGND VPWR VPWR _4946_/X sky130_fd_sc_hd__o2bb2a_1
X_7665_ _7665_/A _7665_/B VGND VGND VPWR VPWR _7682_/A sky130_fd_sc_hd__nor2_1
X_4877_ _4643_/A _4856_/B _4608_/B VGND VGND VPWR VPWR _4877_/Y sky130_fd_sc_hd__a21oi_1
X_7596_ _7475_/X _7522_/B _7593_/X _7594_/Y VGND VGND VPWR VPWR _7686_/A sky130_fd_sc_hd__a211oi_2
X_6616_ _6616_/A _6616_/B _6616_/C VGND VGND VPWR VPWR _6716_/B sky130_fd_sc_hd__and3_1
X_6547_ _6546_/A _6546_/B _6546_/C VGND VGND VPWR VPWR _6548_/C sky130_fd_sc_hd__a21oi_2
X_6478_ _6478_/A _6478_/B VGND VGND VPWR VPWR _6479_/A sky130_fd_sc_hd__and2_1
X_8217_ _8217_/A _8217_/B _8216_/Y VGND VGND VPWR VPWR _8219_/A sky130_fd_sc_hd__nor3b_1
X_5429_ _5364_/X _5428_/X _5481_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
X_9197_ _9224_/CLK _9197_/D VGND VGND VPWR VPWR _9197_/Q sky130_fd_sc_hd__dfxtp_4
X_8148_ _8148_/A VGND VGND VPWR VPWR _8542_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8079_ _8164_/A _8079_/B VGND VGND VPWR VPWR _8081_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4800_ _5738_/S VGND VGND VPWR VPWR _5671_/S sky130_fd_sc_hd__buf_2
XFILLER_34_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5780_ _4608_/B _5713_/S _4608_/X _5779_/X _5676_/A VGND VGND VPWR VPWR _5780_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4731_ _4705_/A _4727_/X _4834_/A VGND VGND VPWR VPWR _4731_/X sky130_fd_sc_hd__mux2_1
X_7450_ _7447_/X _7559_/A _7317_/B _7449_/X VGND VGND VPWR VPWR _7527_/A sky130_fd_sc_hd__o211a_1
X_4662_ _9098_/Q VGND VGND VPWR VPWR _4789_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6401_ _9204_/Q VGND VGND VPWR VPWR _7462_/A sky130_fd_sc_hd__buf_2
X_7381_ _7380_/A _7416_/A _7378_/Y _7379_/X VGND VGND VPWR VPWR _7382_/B sky130_fd_sc_hd__a2bb2o_1
X_9120_ _9216_/CLK hold19/X VGND VGND VPWR VPWR _9120_/Q sky130_fd_sc_hd__dfxtp_2
X_4593_ _4593_/A VGND VGND VPWR VPWR _5432_/A sky130_fd_sc_hd__buf_2
X_6332_ _6332_/A _6332_/B _6332_/C VGND VGND VPWR VPWR _6347_/B sky130_fd_sc_hd__nand3_1
XFILLER_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9051_ _9049_/A _9049_/B _9050_/X VGND VGND VPWR VPWR _9112_/D sky130_fd_sc_hd__a21bo_1
X_6263_ _6263_/A _6263_/B _6263_/C VGND VGND VPWR VPWR _6263_/X sky130_fd_sc_hd__and3_1
X_8002_ _8002_/A _8002_/B VGND VGND VPWR VPWR _8003_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5214_ _5214_/A VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6194_ _6359_/A VGND VGND VPWR VPWR _6968_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5145_ _5656_/B VGND VGND VPWR VPWR _5369_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _4963_/A _5080_/C _5080_/B VGND VGND VPWR VPWR _5076_/X sky130_fd_sc_hd__o21ba_1
X_8904_ _8904_/A _8904_/B _8904_/C VGND VGND VPWR VPWR _8905_/B sky130_fd_sc_hd__and3_1
XFILLER_25_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8835_ _8836_/A _8836_/B _8836_/C VGND VGND VPWR VPWR _8889_/A sky130_fd_sc_hd__o21ai_1
XFILLER_25_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8766_ _8776_/A _8776_/B VGND VGND VPWR VPWR _8766_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5978_ _5915_/A _5915_/C _5915_/B VGND VGND VPWR VPWR _5979_/C sky130_fd_sc_hd__a21bo_1
X_8697_ _8624_/X _8697_/B _8697_/C VGND VGND VPWR VPWR _8699_/A sky130_fd_sc_hd__and3b_1
X_7717_ _7718_/A _7718_/B VGND VGND VPWR VPWR _7717_/X sky130_fd_sc_hd__and2_1
X_4929_ _4929_/A _4929_/B VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7648_ _7770_/A _7769_/A VGND VGND VPWR VPWR _7648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7579_ _8052_/B VGND VGND VPWR VPWR _8467_/A sky130_fd_sc_hd__buf_2
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6950_ _6959_/A _6959_/B VGND VGND VPWR VPWR _6957_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5901_ _9194_/Q _9167_/Q VGND VGND VPWR VPWR _5903_/A sky130_fd_sc_hd__and2_1
X_6881_ _6882_/A _6882_/B _6882_/C _6960_/A VGND VGND VPWR VPWR _6944_/A sky130_fd_sc_hd__o22a_1
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8620_ _8620_/A _8620_/B VGND VGND VPWR VPWR _8622_/B sky130_fd_sc_hd__nand2_1
X_5832_ _5832_/A VGND VGND VPWR VPWR _5833_/A sky130_fd_sc_hd__inv_2
X_8551_ _8551_/A _8551_/B VGND VGND VPWR VPWR _8552_/B sky130_fd_sc_hd__or2_1
XFILLER_61_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5763_ _5583_/X _5632_/X _5765_/A _5762_/Y VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7502_ _7988_/B VGND VGND VPWR VPWR _8091_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4714_ _4705_/A _4712_/X _5730_/S VGND VGND VPWR VPWR _4714_/X sky130_fd_sc_hd__mux2_1
X_8482_ _8363_/A _8482_/B VGND VGND VPWR VPWR _8482_/X sky130_fd_sc_hd__and2b_1
X_5694_ _4643_/A _5693_/X _5738_/S VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__mux2_1
X_7433_ _7822_/D VGND VGND VPWR VPWR _8050_/D sky130_fd_sc_hd__clkbuf_2
X_4645_ _9094_/Q VGND VGND VPWR VPWR _4783_/A sky130_fd_sc_hd__clkbuf_2
X_7364_ _9183_/Q VGND VGND VPWR VPWR _7986_/B sky130_fd_sc_hd__clkbuf_2
X_4576_ _9092_/Q VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__clkbuf_2
X_6315_ _7325_/A VGND VGND VPWR VPWR _7808_/B sky130_fd_sc_hd__buf_2
X_9103_ _9116_/CLK _9103_/D VGND VGND VPWR VPWR _9103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9034_ _9041_/A _9041_/B VGND VGND VPWR VPWR _9035_/C sky130_fd_sc_hd__xnor2_1
X_7295_ _7293_/X _9213_/Q _7295_/C _7295_/D VGND VGND VPWR VPWR _7296_/B sky130_fd_sc_hd__and4b_1
XFILLER_103_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6246_ _6163_/A _6163_/B _6163_/C VGND VGND VPWR VPWR _6248_/C sky130_fd_sc_hd__a21bo_1
XFILLER_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6177_ _9201_/Q VGND VGND VPWR VPWR _6607_/B sky130_fd_sc_hd__buf_2
X_5128_ _5211_/A VGND VGND VPWR VPWR _5630_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5059_ _5621_/A _5055_/X _5057_/X _5258_/A VGND VGND VPWR VPWR _5059_/X sky130_fd_sc_hd__a211o_1
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8818_ _8830_/A _8818_/B VGND VGND VPWR VPWR _8819_/C sky130_fd_sc_hd__xnor2_1
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8749_ _8778_/A _8749_/B VGND VGND VPWR VPWR _8777_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X VGND VGND VPWR VPWR _9216_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA_2 _9191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6100_ _6100_/A _6100_/B VGND VGND VPWR VPWR _6101_/B sky130_fd_sc_hd__xnor2_1
X_7080_ _7039_/A _7038_/A _7038_/B VGND VGND VPWR VPWR _7086_/A sky130_fd_sc_hd__o21ba_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6031_ _6031_/A _7129_/A VGND VGND VPWR VPWR _6032_/B sky130_fd_sc_hd__nand2_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7982_ _8239_/D VGND VGND VPWR VPWR _8717_/A sky130_fd_sc_hd__buf_2
XFILLER_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6933_ _6933_/A _6933_/B VGND VGND VPWR VPWR _6934_/C sky130_fd_sc_hd__xnor2_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6864_ _6864_/A _6864_/B VGND VGND VPWR VPWR _6868_/A sky130_fd_sc_hd__xnor2_1
X_8603_ _8603_/A _8603_/B VGND VGND VPWR VPWR _8604_/B sky130_fd_sc_hd__and2_1
X_5815_ _6022_/A VGND VGND VPWR VPWR _6859_/B sky130_fd_sc_hd__clkbuf_2
X_6795_ _6795_/A _6795_/B _6795_/C VGND VGND VPWR VPWR _6808_/B sky130_fd_sc_hd__nand3_1
X_8534_ _8451_/A _8456_/B _8451_/B VGND VGND VPWR VPWR _8535_/B sky130_fd_sc_hd__o21ba_1
X_5746_ _5424_/X _5558_/X _5420_/X _4676_/C VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__o22a_1
XFILLER_41_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8465_ _8465_/A _8465_/B VGND VGND VPWR VPWR _8469_/A sky130_fd_sc_hd__nor2_1
X_5677_ _5124_/X _4812_/X _5204_/A _5675_/X _5676_/Y VGND VGND VPWR VPWR _9146_/D
+ sky130_fd_sc_hd__o221a_1
X_7416_ _7416_/A VGND VGND VPWR VPWR _7447_/B sky130_fd_sc_hd__clkinv_2
X_4628_ _4799_/A VGND VGND VPWR VPWR _4629_/A sky130_fd_sc_hd__buf_2
X_8396_ _8397_/A _8397_/B VGND VGND VPWR VPWR _8396_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7347_ _7347_/A _7347_/B VGND VGND VPWR VPWR _7347_/Y sky130_fd_sc_hd__nand2_1
X_4559_ _4874_/S VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7278_ _7276_/X _7277_/Y _7168_/Y _7171_/B VGND VGND VPWR VPWR _7284_/B sky130_fd_sc_hd__o211ai_1
X_9017_ _9017_/A _9023_/A VGND VGND VPWR VPWR _9038_/A sky130_fd_sc_hd__xnor2_2
X_6229_ _6145_/A _6145_/C _6145_/B VGND VGND VPWR VPWR _6231_/C sky130_fd_sc_hd__a21bo_1
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR clkbuf_4_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
Xoutput94 _9136_/Q VGND VGND VPWR VPWR F[7] sky130_fd_sc_hd__buf_2
Xoutput83 _9155_/Q VGND VGND VPWR VPWR F[26] sky130_fd_sc_hd__buf_2
Xoutput72 _9145_/Q VGND VGND VPWR VPWR F[16] sky130_fd_sc_hd__buf_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5600_ _5484_/A _5599_/X _5695_/S VGND VGND VPWR VPWR _5600_/X sky130_fd_sc_hd__mux2_1
X_6580_ _6580_/A _6580_/B _6580_/C VGND VGND VPWR VPWR _6582_/A sky130_fd_sc_hd__nand3_1
X_5531_ _5484_/X _5530_/X _5603_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
X_8250_ _8157_/A _8159_/B _8157_/B VGND VGND VPWR VPWR _8361_/A sky130_fd_sc_hd__o21ba_1
X_7201_ _7201_/A _7309_/B VGND VGND VPWR VPWR _7202_/B sky130_fd_sc_hd__nand2_1
X_5462_ _9078_/Q _5559_/B VGND VGND VPWR VPWR _5462_/Y sky130_fd_sc_hd__nor2_1
X_8181_ _8316_/B _8181_/B VGND VGND VPWR VPWR _8183_/A sky130_fd_sc_hd__xnor2_1
X_5393_ _5393_/A VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__inv_2
X_7132_ _7132_/A _7132_/B VGND VGND VPWR VPWR _7133_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7063_ _7072_/A _7072_/B VGND VGND VPWR VPWR _7064_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6014_ _6014_/A VGND VGND VPWR VPWR _6859_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7965_ _6192_/X _8150_/D _8607_/C _8156_/A VGND VGND VPWR VPWR _7967_/A sky130_fd_sc_hd__a22oi_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7896_ _7779_/A _7779_/B _7895_/Y VGND VGND VPWR VPWR _8009_/B sky130_fd_sc_hd__a21o_2
X_6916_ _6808_/C _6809_/B _6912_/Y _6914_/Y VGND VGND VPWR VPWR _7054_/A sky130_fd_sc_hd__a211oi_4
X_6847_ _6847_/A _6850_/B VGND VGND VPWR VPWR _6848_/B sky130_fd_sc_hd__xor2_2
X_6778_ _6886_/A _6778_/B _7465_/A _7360_/A VGND VGND VPWR VPWR _6780_/A sky130_fd_sc_hd__and4_1
X_8517_ _8517_/A _8664_/D _8660_/C VGND VGND VPWR VPWR _8518_/B sky130_fd_sc_hd__and3_1
X_5729_ _4582_/A _5728_/X _5729_/S VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8448_ _8556_/A _8448_/B VGND VGND VPWR VPWR _8487_/A sky130_fd_sc_hd__or2_1
X_8379_ _8379_/A VGND VGND VPWR VPWR _8527_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7750_ _8464_/B VGND VGND VPWR VPWR _8677_/A sky130_fd_sc_hd__buf_2
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4962_ _4642_/A _4959_/X _4960_/X _4961_/X VGND VGND VPWR VPWR _4962_/X sky130_fd_sc_hd__o22a_1
X_7681_ _7562_/A _8639_/B _7563_/A _7561_/B VGND VGND VPWR VPWR _7791_/A sky130_fd_sc_hd__a31o_1
X_6701_ _6701_/A _6701_/B VGND VGND VPWR VPWR _6709_/A sky130_fd_sc_hd__xnor2_2
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4893_ _5282_/S _4856_/B _4892_/X VGND VGND VPWR VPWR _4893_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6632_ _7389_/A _8780_/A _6632_/C VGND VGND VPWR VPWR _6734_/A sky130_fd_sc_hd__and3_1
X_6563_ _6506_/B _6563_/B VGND VGND VPWR VPWR _6563_/X sky130_fd_sc_hd__and2b_1
X_8302_ _8196_/A _8196_/B _8301_/X VGND VGND VPWR VPWR _8304_/B sky130_fd_sc_hd__a21oi_1
X_5514_ _4847_/A _5211_/A _5513_/X _4584_/A VGND VGND VPWR VPWR _5514_/Y sky130_fd_sc_hd__a211oi_1
X_6494_ _7187_/B _6493_/C _7604_/D _6858_/A VGND VGND VPWR VPWR _6495_/B sky130_fd_sc_hd__a22o_1
X_8233_ _8226_/A _8233_/B VGND VGND VPWR VPWR _8331_/A sky130_fd_sc_hd__and2b_1
X_5445_ _5385_/X _5389_/X _4656_/A VGND VGND VPWR VPWR _5445_/Y sky130_fd_sc_hd__a21oi_1
X_8164_ _8164_/A _8164_/B VGND VGND VPWR VPWR _8165_/B sky130_fd_sc_hd__or2_2
X_7115_ _7499_/A _7610_/D _7246_/A _7114_/Y VGND VGND VPWR VPWR _7117_/A sky130_fd_sc_hd__o2bb2a_1
X_5376_ _5249_/X _5246_/Y _5258_/X VGND VGND VPWR VPWR _5376_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8095_ _7967_/A _7970_/B _7967_/B VGND VGND VPWR VPWR _8096_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7046_ _7143_/B _7046_/B VGND VGND VPWR VPWR _7047_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8997_ _8958_/B _8973_/X _8995_/Y _8996_/X VGND VGND VPWR VPWR _8999_/A sky130_fd_sc_hd__o211a_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _7948_/A _7948_/B VGND VGND VPWR VPWR _7950_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7879_ _7770_/C _7771_/A _7648_/Y VGND VGND VPWR VPWR _7887_/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5230_ _9104_/Q VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5161_ _9075_/Q VGND VGND VPWR VPWR _5370_/A sky130_fd_sc_hd__clkinv_2
X_5092_ _5087_/X _5088_/Y _5089_/X _5090_/X _5091_/Y VGND VGND VPWR VPWR _5092_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8920_ _8920_/A _8920_/B VGND VGND VPWR VPWR _8965_/A sky130_fd_sc_hd__xnor2_1
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8851_ _8852_/A _8852_/B VGND VGND VPWR VPWR _8853_/A sky130_fd_sc_hd__or2_1
XFILLER_64_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8782_ _8782_/A _8842_/B VGND VGND VPWR VPWR _8784_/B sky130_fd_sc_hd__and2_1
X_7802_ _7801_/A _7801_/B _7800_/Y VGND VGND VPWR VPWR _7803_/B sky130_fd_sc_hd__o21ba_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5994_ _6037_/A _6037_/C _6037_/B VGND VGND VPWR VPWR _5994_/Y sky130_fd_sc_hd__a21oi_1
X_7733_ _8091_/A _8091_/B _7959_/D _7748_/A VGND VGND VPWR VPWR _7734_/B sky130_fd_sc_hd__and4_1
X_4945_ _4934_/X _4941_/X _4944_/Y _4570_/A _5007_/A VGND VGND VPWR VPWR _4945_/X
+ sky130_fd_sc_hd__o221a_1
X_7664_ _7691_/A _7691_/B VGND VGND VPWR VPWR _7666_/A sky130_fd_sc_hd__xor2_1
X_4876_ _4876_/A _4876_/B VGND VGND VPWR VPWR _4876_/Y sky130_fd_sc_hd__nand2_1
X_7595_ _7593_/X _7594_/Y _7475_/X _7522_/B VGND VGND VPWR VPWR _7684_/B sky130_fd_sc_hd__o211ai_1
X_6615_ _6615_/A _6691_/B VGND VGND VPWR VPWR _6616_/C sky130_fd_sc_hd__nand2_1
XFILLER_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6546_ _6546_/A _6546_/B _6546_/C VGND VGND VPWR VPWR _6548_/B sky130_fd_sc_hd__and3_1
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6477_ _6476_/A _6476_/B _6476_/C VGND VGND VPWR VPWR _6478_/B sky130_fd_sc_hd__o21ai_1
X_8216_ _8220_/A _8933_/B _8045_/A _8215_/X VGND VGND VPWR VPWR _8216_/Y sky130_fd_sc_hd__a31oi_1
X_5428_ _5339_/X _5427_/X _5428_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
X_9196_ _9216_/CLK _9196_/D VGND VGND VPWR VPWR _9196_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8147_ _8516_/A VGND VGND VPWR VPWR _8337_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5359_ _5628_/A VGND VGND VPWR VPWR _5481_/S sky130_fd_sc_hd__clkbuf_2
X_8078_ _8078_/A _8078_/B _8078_/C VGND VGND VPWR VPWR _8079_/B sky130_fd_sc_hd__or3_1
XFILLER_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7029_ _7029_/A _7029_/B _7029_/C VGND VGND VPWR VPWR _7053_/B sky130_fd_sc_hd__and3_2
XFILLER_74_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4730_ _5692_/S VGND VGND VPWR VPWR _4834_/A sky130_fd_sc_hd__clkbuf_2
X_4661_ _4661_/A VGND VGND VPWR VPWR _5364_/A sky130_fd_sc_hd__clkbuf_2
X_7380_ _7380_/A _7416_/A _7378_/Y _7379_/X VGND VGND VPWR VPWR _7382_/A sky130_fd_sc_hd__or4bb_2
X_6400_ _6825_/A VGND VGND VPWR VPWR _7295_/C sky130_fd_sc_hd__clkbuf_2
X_4592_ _5156_/A VGND VGND VPWR VPWR _4593_/A sky130_fd_sc_hd__clkbuf_2
X_6331_ _6434_/A _6434_/B VGND VGND VPWR VPWR _6332_/C sky130_fd_sc_hd__xnor2_1
X_9050_ _9046_/A _9045_/B _9045_/A VGND VGND VPWR VPWR _9050_/X sky130_fd_sc_hd__o21ba_1
XFILLER_6_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6262_ _6263_/B _6263_/C _6263_/A VGND VGND VPWR VPWR _6262_/Y sky130_fd_sc_hd__a21oi_1
X_8001_ _8001_/A _8001_/B VGND VGND VPWR VPWR _8002_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5213_ _5213_/A VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6193_ _7299_/A _8349_/A _6192_/X _6358_/A VGND VGND VPWR VPWR _6202_/A sky130_fd_sc_hd__a22oi_2
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5144_ _5144_/A VGND VGND VPWR VPWR _5313_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5075_ _5169_/A _5073_/Y _5074_/X _4548_/A VGND VGND VPWR VPWR _5075_/X sky130_fd_sc_hd__a31o_1
X_8903_ _8904_/A _8904_/B _8904_/C VGND VGND VPWR VPWR _8947_/A sky130_fd_sc_hd__a21oi_1
XFILLER_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8834_ _8937_/A _8937_/B _8833_/X VGND VGND VPWR VPWR _8836_/C sky130_fd_sc_hd__o21a_1
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8765_ _8700_/A _8989_/B _8701_/A _8699_/B VGND VGND VPWR VPWR _8776_/B sky130_fd_sc_hd__a31o_1
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5977_ _5976_/A _5976_/C _5976_/B VGND VGND VPWR VPWR _5979_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8696_ _8600_/A _8600_/B _8604_/B VGND VGND VPWR VPWR _8697_/C sky130_fd_sc_hd__a21oi_1
X_7716_ _7716_/A _7716_/B VGND VGND VPWR VPWR _7718_/B sky130_fd_sc_hd__xnor2_1
X_4928_ _4928_/A _4939_/B VGND VGND VPWR VPWR _4929_/B sky130_fd_sc_hd__nand2_1
X_7647_ _7647_/A _8243_/B VGND VGND VPWR VPWR _7770_/C sky130_fd_sc_hd__nand2_1
XFILLER_60_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4859_ _4847_/X _4855_/X _4856_/Y _5251_/A VGND VGND VPWR VPWR _4859_/X sky130_fd_sc_hd__o211a_1
X_7578_ _7810_/C VGND VGND VPWR VPWR _8032_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6529_ _6590_/B _7706_/B _6886_/B _7016_/A VGND VGND VPWR VPWR _6531_/A sky130_fd_sc_hd__a22oi_2
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9179_ _9213_/CLK input9/X VGND VGND VPWR VPWR _9179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _9165_/Q _6447_/A _6055_/A _9166_/Q VGND VGND VPWR VPWR _5903_/C sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _6879_/A _6940_/B _6879_/C VGND VGND VPWR VPWR _6960_/A sky130_fd_sc_hd__o21a_1
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5831_ _7293_/B _6151_/A _6590_/B _6031_/A VGND VGND VPWR VPWR _5832_/A sky130_fd_sc_hd__a22o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8550_ _8551_/A _8551_/B VGND VGND VPWR VPWR _8552_/A sky130_fd_sc_hd__nand2_1
X_5762_ _4876_/A _5606_/X _5632_/A VGND VGND VPWR VPWR _5762_/Y sky130_fd_sc_hd__a21oi_1
X_7501_ _7880_/A _7966_/D VGND VGND VPWR VPWR _7501_/Y sky130_fd_sc_hd__nand2_1
X_4713_ _9099_/Q VGND VGND VPWR VPWR _5730_/S sky130_fd_sc_hd__inv_2
X_8481_ _8481_/A _8481_/B VGND VGND VPWR VPWR _8481_/Y sky130_fd_sc_hd__nor2_1
X_5693_ _4637_/A _5692_/X _5737_/S VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7432_ _7329_/A _7328_/A _7328_/B VGND VGND VPWR VPWR _7439_/A sky130_fd_sc_hd__o21ba_1
X_4644_ _5402_/A _5484_/A _5534_/A _5557_/A VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__or4_1
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7363_ _7482_/B _7363_/B VGND VGND VPWR VPWR _7496_/A sky130_fd_sc_hd__nor2_1
X_4575_ _4780_/A VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__inv_2
X_6314_ _6760_/A VGND VGND VPWR VPWR _7325_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9102_ _9223_/CLK _9102_/D VGND VGND VPWR VPWR _9102_/Q sky130_fd_sc_hd__dfxtp_1
X_7294_ _7295_/C _9213_/Q _7292_/Y _7293_/X VGND VGND VPWR VPWR _7296_/A sky130_fd_sc_hd__o2bb2a_1
X_9033_ _9006_/A _9006_/B _9008_/A _9008_/B VGND VGND VPWR VPWR _9041_/B sky130_fd_sc_hd__o22a_1
X_6245_ _6245_/A _6245_/B _6332_/A VGND VGND VPWR VPWR _6332_/B sky130_fd_sc_hd__nand3_2
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6176_ _6825_/A VGND VGND VPWR VPWR _6567_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5127_ _9082_/Q VGND VGND VPWR VPWR _5211_/A sky130_fd_sc_hd__buf_2
X_5058_ _5058_/A VGND VGND VPWR VPWR _5258_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8817_ _8817_/A _8817_/B VGND VGND VPWR VPWR _8818_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8748_ _8814_/A _8778_/C VGND VGND VPWR VPWR _8749_/B sky130_fd_sc_hd__nor2_1
XFILLER_71_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8679_ _8816_/A _8794_/B VGND VGND VPWR VPWR _8680_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _9191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6030_ _9201_/Q VGND VGND VPWR VPWR _7129_/A sky130_fd_sc_hd__clkbuf_2
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7981_ _7981_/A _8064_/B VGND VGND VPWR VPWR _8003_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6932_ _7031_/B _6932_/B VGND VGND VPWR VPWR _6933_/B sky130_fd_sc_hd__xnor2_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6863_ _6982_/A _6863_/B VGND VGND VPWR VPWR _6864_/B sky130_fd_sc_hd__xnor2_1
X_8602_ _8603_/A _8603_/B VGND VGND VPWR VPWR _8604_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5814_ _9164_/Q VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__clkbuf_2
X_6794_ _6884_/A _6884_/B VGND VGND VPWR VPWR _6795_/C sky130_fd_sc_hd__xnor2_1
X_8533_ _8533_/A _8533_/B VGND VGND VPWR VPWR _8633_/B sky130_fd_sc_hd__nor2_1
X_5745_ _5745_/A VGND VGND VPWR VPWR _9149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8464_ _8664_/A _8464_/B _8664_/B _8674_/A VGND VGND VPWR VPWR _8465_/B sky130_fd_sc_hd__and4_1
X_5676_ _5676_/A _5676_/B VGND VGND VPWR VPWR _5676_/Y sky130_fd_sc_hd__nand2_1
X_7415_ _7340_/A _7340_/B _7340_/C VGND VGND VPWR VPWR _7447_/A sky130_fd_sc_hd__a21o_2
X_4627_ _9106_/Q VGND VGND VPWR VPWR _4799_/A sky130_fd_sc_hd__clkbuf_2
X_8395_ _8395_/A _8395_/B VGND VGND VPWR VPWR _8397_/B sky130_fd_sc_hd__nand2_1
X_7346_ _9201_/Q _7346_/B VGND VGND VPWR VPWR _7351_/A sky130_fd_sc_hd__nand2_1
X_4558_ _4558_/A VGND VGND VPWR VPWR _4874_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7277_ _7277_/A _7394_/B _7277_/C _7277_/D VGND VGND VPWR VPWR _7277_/Y sky130_fd_sc_hd__nor4_4
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9016_ _8989_/A _8989_/B _8990_/A _9015_/X VGND VGND VPWR VPWR _9023_/A sky130_fd_sc_hd__a31oi_4
X_6228_ _7509_/A _7602_/A _6329_/A _6228_/D VGND VGND VPWR VPWR _6329_/B sky130_fd_sc_hd__nand4_4
X_6159_ _7254_/C VGND VGND VPWR VPWR _6775_/A sky130_fd_sc_hd__buf_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput73 _9146_/Q VGND VGND VPWR VPWR F[17] sky130_fd_sc_hd__buf_2
Xoutput84 _9156_/Q VGND VGND VPWR VPWR F[27] sky130_fd_sc_hd__buf_2
Xoutput95 _9137_/Q VGND VGND VPWR VPWR F[8] sky130_fd_sc_hd__buf_2
XFILLER_76_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5530_ _5461_/X _5529_/X _5553_/S VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
X_5461_ _5749_/A VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7200_ _7200_/A _7200_/B VGND VGND VPWR VPWR _7202_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8180_ _8037_/A _8041_/B _8037_/B VGND VGND VPWR VPWR _8181_/B sky130_fd_sc_hd__o21ba_1
X_5392_ _4883_/X _5117_/A _5387_/X _5390_/Y _5391_/X VGND VGND VPWR VPWR _5392_/X
+ sky130_fd_sc_hd__a221o_1
X_7131_ _7131_/A _7347_/A _7131_/C _7131_/D VGND VGND VPWR VPWR _7132_/B sky130_fd_sc_hd__and4_1
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7062_ _6949_/A _6948_/A _6948_/B VGND VGND VPWR VPWR _7072_/B sky130_fd_sc_hd__o21ba_2
X_6013_ _6013_/A _6013_/B VGND VGND VPWR VPWR _6016_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7964_ _7966_/D VGND VGND VPWR VPWR _8607_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_94_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6915_ _6912_/Y _6914_/Y _6808_/C _6809_/B VGND VGND VPWR VPWR _6939_/B sky130_fd_sc_hd__o211a_1
X_7895_ _7895_/A _7895_/B VGND VGND VPWR VPWR _7895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6846_ _6744_/A _6744_/B _6845_/X VGND VGND VPWR VPWR _6850_/B sky130_fd_sc_hd__o21bai_2
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6777_ _7119_/C VGND VGND VPWR VPWR _7360_/A sky130_fd_sc_hd__buf_2
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8516_ _8516_/A _8516_/B VGND VGND VPWR VPWR _8660_/C sky130_fd_sc_hd__and2_1
XFILLER_50_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5728_ _9094_/Q _5727_/X _5728_/S VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__mux2_1
X_8447_ _8447_/A _8447_/B _8447_/C VGND VGND VPWR VPWR _8448_/B sky130_fd_sc_hd__nor3_1
X_5659_ _4584_/A _5420_/A _4861_/A VGND VGND VPWR VPWR _5659_/Y sky130_fd_sc_hd__a21oi_1
X_8378_ _8297_/A _8378_/B VGND VGND VPWR VPWR _8393_/A sky130_fd_sc_hd__and2b_1
X_7329_ _7329_/A _7329_/B VGND VGND VPWR VPWR _7338_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X VGND VGND VPWR VPWR _9213_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_92_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4961_ _4827_/B _4957_/B _5733_/S VGND VGND VPWR VPWR _4961_/X sky130_fd_sc_hd__a21o_1
X_7680_ _8816_/B VGND VGND VPWR VPWR _8639_/B sky130_fd_sc_hd__buf_2
X_6700_ _6700_/A _7849_/B VGND VGND VPWR VPWR _6701_/B sky130_fd_sc_hd__nand2_1
X_4892_ _4538_/A _4830_/X _4888_/X _4890_/Y _4891_/X VGND VGND VPWR VPWR _4892_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6631_ _7194_/A _8584_/A _6495_/B _6493_/X VGND VGND VPWR VPWR _6632_/C sky130_fd_sc_hd__a31o_1
X_8301_ _8195_/A _8301_/B VGND VGND VPWR VPWR _8301_/X sky130_fd_sc_hd__and2b_1
X_6562_ _6649_/A _6562_/B VGND VGND VPWR VPWR _9081_/D sky130_fd_sc_hd__nor2_1
X_5513_ _5131_/A _4579_/A _4659_/A _9079_/Q _5512_/Y VGND VGND VPWR VPWR _5513_/X
+ sky130_fd_sc_hd__o221a_1
X_6493_ _7187_/B _7093_/B _6493_/C _7604_/D VGND VGND VPWR VPWR _6493_/X sky130_fd_sc_hd__and4_1
X_8232_ _8232_/A _8232_/B VGND VGND VPWR VPWR _9096_/D sky130_fd_sc_hd__xnor2_1
X_5444_ _5266_/X _5206_/A _5442_/X _5443_/Y _4550_/A VGND VGND VPWR VPWR _5444_/X
+ sky130_fd_sc_hd__a221o_1
X_8163_ _8164_/A _8164_/B VGND VGND VPWR VPWR _8165_/A sky130_fd_sc_hd__nand2_1
X_7114_ _5908_/B _7348_/B _7640_/A _6240_/A VGND VGND VPWR VPWR _7114_/Y sky130_fd_sc_hd__a22oi_1
X_5375_ _5368_/X _5555_/A _5373_/X _5374_/Y _4593_/A VGND VGND VPWR VPWR _5375_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8094_ _8094_/A _8094_/B VGND VGND VPWR VPWR _8146_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7045_ _6930_/A _6929_/B _6929_/A VGND VGND VPWR VPWR _7046_/B sky130_fd_sc_hd__o21ba_1
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8996_ _8948_/A _8952_/B _8993_/X _9018_/A VGND VGND VPWR VPWR _8996_/X sky130_fd_sc_hd__a211o_1
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A VGND VGND VPWR VPWR clkbuf_4_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_7947_ _7946_/A _7946_/B _7945_/X VGND VGND VPWR VPWR _7948_/B sky130_fd_sc_hd__o21bai_2
X_7878_ _7878_/A _7957_/A VGND VGND VPWR VPWR _7890_/A sky130_fd_sc_hd__xor2_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6829_ _6829_/A _6829_/B VGND VGND VPWR VPWR _6830_/B sky130_fd_sc_hd__xnor2_4
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5160_ _5160_/A VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _4940_/C _4998_/A _5041_/A VGND VGND VPWR VPWR _5091_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8850_ _8909_/A _8850_/B VGND VGND VPWR VPWR _8852_/B sky130_fd_sc_hd__and2_1
X_8781_ _8781_/A _8836_/A VGND VGND VPWR VPWR _8784_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7801_ _7801_/A _7801_/B _7800_/Y VGND VGND VPWR VPWR _7803_/A sky130_fd_sc_hd__nor3b_1
X_5993_ _6037_/A _6037_/B _6037_/C VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__and3_1
X_7732_ _8156_/B _7959_/D _7748_/A _8154_/A VGND VGND VPWR VPWR _7734_/A sky130_fd_sc_hd__a22oi_1
X_4944_ _4944_/A _5093_/A VGND VGND VPWR VPWR _4944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7663_ _7663_/A _7784_/A VGND VGND VPWR VPWR _7691_/B sky130_fd_sc_hd__or2_2
X_4875_ _4830_/X _4874_/X _4875_/S VGND VGND VPWR VPWR _4876_/B sky130_fd_sc_hd__mux2_1
X_7594_ _7594_/A _7594_/B VGND VGND VPWR VPWR _7594_/Y sky130_fd_sc_hd__nor2_1
X_6614_ _6614_/A _6614_/B _6691_/A VGND VGND VPWR VPWR _6691_/B sky130_fd_sc_hd__nand3_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6545_ _6616_/B _6545_/B VGND VGND VPWR VPWR _6546_/C sky130_fd_sc_hd__nand2_2
X_8215_ _8043_/B _8215_/B VGND VGND VPWR VPWR _8215_/X sky130_fd_sc_hd__and2b_1
X_6476_ _6476_/A _6476_/B _6476_/C VGND VGND VPWR VPWR _6478_/A sky130_fd_sc_hd__or3_1
X_5427_ _5315_/X _5426_/X _5427_/S VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__mux2_1
X_9195_ _9220_/CLK _9195_/D VGND VGND VPWR VPWR _9195_/Q sky130_fd_sc_hd__dfxtp_2
X_8146_ _8096_/B _8146_/B VGND VGND VPWR VPWR _8166_/A sky130_fd_sc_hd__and2b_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _5287_/X _5357_/X _5428_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
X_8077_ _8078_/A _8078_/B _8078_/C VGND VGND VPWR VPWR _8164_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7028_ _7028_/A _7141_/B VGND VGND VPWR VPWR _7029_/C sky130_fd_sc_hd__nand2_1
XFILLER_59_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5289_ _5252_/A _9073_/Q _4659_/A _9071_/Q _4571_/A VGND VGND VPWR VPWR _5289_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8979_ _8979_/A _8979_/B VGND VGND VPWR VPWR _8980_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4660_ _4660_/A VGND VGND VPWR VPWR _4676_/C sky130_fd_sc_hd__buf_2
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6330_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6434_/B sky130_fd_sc_hd__xor2_1
X_4591_ _4591_/A VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6261_ _6261_/A _6352_/B VGND VGND VPWR VPWR _6263_/A sky130_fd_sc_hd__xnor2_1
X_8000_ _8001_/A _8001_/B VGND VGND VPWR VPWR _8002_/A sky130_fd_sc_hd__and2_1
XFILLER_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6192_ _8091_/B VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__buf_4
XFILLER_69_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5212_ _5212_/A VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__buf_2
X_5143_ _9072_/Q VGND VGND VPWR VPWR _5362_/A sky130_fd_sc_hd__buf_2
XFILLER_56_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5074_ _5074_/A _5074_/B _5080_/C VGND VGND VPWR VPWR _5074_/X sky130_fd_sc_hd__or3_1
XFILLER_84_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8902_ _8902_/A _8902_/B VGND VGND VPWR VPWR _8904_/C sky130_fd_sc_hd__xnor2_1
X_8833_ _8666_/A _8831_/B _8832_/B _8831_/A VGND VGND VPWR VPWR _8833_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8764_ _9025_/B VGND VGND VPWR VPWR _8989_/B sky130_fd_sc_hd__clkbuf_2
X_5976_ _5976_/A _5976_/B _5976_/C VGND VGND VPWR VPWR _5979_/A sky130_fd_sc_hd__nand3_1
X_8695_ _8695_/A _8761_/A VGND VGND VPWR VPWR _8703_/A sky130_fd_sc_hd__or2_1
X_7715_ _7589_/A _7589_/B _7714_/X VGND VGND VPWR VPWR _7716_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4927_ _4927_/A _5044_/A VGND VGND VPWR VPWR _4980_/B sky130_fd_sc_hd__or2_2
X_7646_ _7986_/B VGND VGND VPWR VPWR _8243_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4858_ _5007_/A VGND VGND VPWR VPWR _5251_/A sky130_fd_sc_hd__clkbuf_2
X_7577_ _7577_/A _7577_/B VGND VGND VPWR VPWR _7594_/A sky130_fd_sc_hd__or2_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4789_ _4789_/A VGND VGND VPWR VPWR _5058_/A sky130_fd_sc_hd__clkbuf_2
X_6528_ _7131_/D VGND VGND VPWR VPWR _6886_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6459_ _6458_/A _6458_/B _6458_/C VGND VGND VPWR VPWR _6546_/A sky130_fd_sc_hd__a21o_1
X_9178_ _9213_/CLK input8/X VGND VGND VPWR VPWR _9178_/Q sky130_fd_sc_hd__dfxtp_1
X_8129_ _8024_/B _8025_/A _8128_/Y _8019_/B _8126_/X VGND VGND VPWR VPWR _8130_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5830_ _6998_/B VGND VGND VPWR VPWR _6590_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5761_ _4889_/X _4535_/X _5756_/X _5760_/X _5765_/B VGND VGND VPWR VPWR _5761_/X
+ sky130_fd_sc_hd__o32a_1
X_7500_ _8091_/C VGND VGND VPWR VPWR _7966_/D sky130_fd_sc_hd__clkbuf_2
X_8480_ _8480_/A _8480_/B VGND VGND VPWR VPWR _8480_/X sky130_fd_sc_hd__or2_2
X_4712_ _4759_/A _4711_/X _5729_/S VGND VGND VPWR VPWR _4712_/X sky130_fd_sc_hd__mux2_1
X_7431_ _7918_/A _8185_/A _7310_/A _7308_/B VGND VGND VPWR VPWR _7440_/A sky130_fd_sc_hd__a31o_1
X_5692_ _5367_/X _5691_/X _5692_/S VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__mux2_1
X_4643_ _4643_/A VGND VGND VPWR VPWR _5557_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7362_ _6775_/A _7756_/A _7358_/Y _7482_/A VGND VGND VPWR VPWR _7363_/B sky130_fd_sc_hd__o2bb2a_1
X_4574_ _9093_/Q VGND VGND VPWR VPWR _4780_/A sky130_fd_sc_hd__clkbuf_2
X_6313_ _6313_/A _6313_/B _6679_/A _7604_/B VGND VGND VPWR VPWR _6320_/A sky130_fd_sc_hd__and4_1
X_9101_ _9223_/CLK _9101_/D VGND VGND VPWR VPWR _9101_/Q sky130_fd_sc_hd__dfxtp_2
X_7293_ _7293_/A _7293_/B _9211_/Q _7419_/D VGND VGND VPWR VPWR _7293_/X sky130_fd_sc_hd__and4_1
X_9032_ _9032_/A _9032_/B VGND VGND VPWR VPWR _9041_/A sky130_fd_sc_hd__xnor2_1
X_6244_ _6245_/B _6332_/A _6245_/A VGND VGND VPWR VPWR _6248_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6175_ _6175_/A _6175_/B VGND VGND VPWR VPWR _6179_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5126_ _5126_/A VGND VGND VPWR VPWR _5126_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5057_ _4845_/Y _5046_/Y _5056_/X _4841_/A VGND VGND VPWR VPWR _5057_/X sky130_fd_sc_hd__o211a_1
XFILLER_72_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8816_ _8816_/A _8816_/B VGND VGND VPWR VPWR _8817_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8747_ _8746_/A _8806_/B _8746_/C VGND VGND VPWR VPWR _8778_/C sky130_fd_sc_hd__a21oi_1
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ _6358_/A VGND VGND VPWR VPWR _7194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8678_ _8678_/A _8678_/B VGND VGND VPWR VPWR _8680_/A sky130_fd_sc_hd__nor2_1
X_7629_ _7629_/A _7629_/B VGND VGND VPWR VPWR _7629_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 _9199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7980_ _7978_/X _7860_/B _7976_/Y _8064_/A VGND VGND VPWR VPWR _8064_/B sky130_fd_sc_hd__o211ai_4
XFILLER_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6931_ _6763_/A _6762_/B _6762_/A VGND VGND VPWR VPWR _6932_/B sky130_fd_sc_hd__o21ba_1
X_6862_ _6862_/A _6862_/B VGND VGND VPWR VPWR _6863_/B sky130_fd_sc_hd__xnor2_1
X_5813_ _7257_/A VGND VGND VPWR VPWR _7509_/A sky130_fd_sc_hd__buf_4
X_8601_ _8700_/A _8798_/B VGND VGND VPWR VPWR _8603_/B sky130_fd_sc_hd__and2_1
XFILLER_62_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8532_ _8530_/X _8846_/B _8700_/A _8532_/D VGND VGND VPWR VPWR _8533_/B sky130_fd_sc_hd__and4b_1
X_6793_ _6793_/A _6883_/A VGND VGND VPWR VPWR _6884_/B sky130_fd_sc_hd__xnor2_1
X_5744_ _5206_/X _5743_/X _5785_/S VGND VGND VPWR VPWR _5745_/A sky130_fd_sc_hd__mux2_1
X_8463_ _8675_/A _8831_/A _8674_/A _8780_/A VGND VGND VPWR VPWR _8465_/A sky130_fd_sc_hd__a22oi_1
X_5675_ _5632_/X _5674_/X _5698_/S VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__mux2_1
X_8394_ _8393_/A _8393_/B _8392_/Y VGND VGND VPWR VPWR _8395_/B sky130_fd_sc_hd__o21bai_2
X_4626_ _9112_/Q VGND VGND VPWR VPWR _4982_/A sky130_fd_sc_hd__inv_2
X_7414_ _7389_/A _8867_/B _7397_/B _7396_/B VGND VGND VPWR VPWR _7543_/A sky130_fd_sc_hd__a31oi_2
X_7345_ _7245_/A _7244_/A _7244_/B VGND VGND VPWR VPWR _7452_/A sky130_fd_sc_hd__o21ba_1
X_4557_ _5378_/A VGND VGND VPWR VPWR _4558_/A sky130_fd_sc_hd__clkbuf_2
X_7276_ _7277_/A _7394_/B _7277_/C _7277_/D VGND VGND VPWR VPWR _7276_/X sky130_fd_sc_hd__o22a_1
X_9015_ _8988_/B _9015_/B VGND VGND VPWR VPWR _9015_/X sky130_fd_sc_hd__and2b_1
X_6227_ _7822_/A VGND VGND VPWR VPWR _7602_/A sky130_fd_sc_hd__buf_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6500_/B VGND VGND VPWR VPWR _7309_/A sky130_fd_sc_hd__buf_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5043_/A _5043_/B _5743_/S VGND VGND VPWR VPWR _5109_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6089_ _6090_/A _6090_/B _6090_/C VGND VGND VPWR VPWR _6104_/B sky130_fd_sc_hd__a21o_1
XFILLER_85_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput74 _9147_/Q VGND VGND VPWR VPWR F[18] sky130_fd_sc_hd__buf_2
Xoutput85 _9157_/Q VGND VGND VPWR VPWR F[28] sky130_fd_sc_hd__buf_2
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput96 _9138_/Q VGND VGND VPWR VPWR F[9] sky130_fd_sc_hd__buf_2
XFILLER_91_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5460_ _5460_/A VGND VGND VPWR VPWR _5749_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5391_ _5391_/A VGND VGND VPWR VPWR _5391_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7130_ _5985_/D _7241_/B _7346_/B _6172_/A VGND VGND VPWR VPWR _7132_/A sky130_fd_sc_hd__a22oi_2
X_7061_ _7061_/A _7061_/B VGND VGND VPWR VPWR _7072_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6012_ _6169_/A _7253_/A _7253_/B _9170_/Q VGND VGND VPWR VPWR _6013_/B sky130_fd_sc_hd__and4_1
.ends

