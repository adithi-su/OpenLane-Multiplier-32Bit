VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MULTI_32bit
  CLASS BLOCK ;
  FOREIGN MULTI_32bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 301.290 BY 312.010 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 308.010 203.230 312.010 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 308.010 290.170 312.010 ;
    END
  END A[12]
  PIN A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 258.440 301.290 259.040 ;
    END
  END A[13]
  PIN A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 193.840 301.290 194.440 ;
    END
  END A[14]
  PIN A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END A[15]
  PIN A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 308.010 106.630 312.010 ;
    END
  END A[16]
  PIN A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 308.010 119.510 312.010 ;
    END
  END A[17]
  PIN A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END A[18]
  PIN A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 299.240 301.290 299.840 ;
    END
  END A[19]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 78.240 301.290 78.840 ;
    END
  END A[1]
  PIN A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 248.240 301.290 248.840 ;
    END
  END A[20]
  PIN A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 308.010 93.750 312.010 ;
    END
  END A[21]
  PIN A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END A[22]
  PIN A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END A[23]
  PIN A[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END A[24]
  PIN A[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 285.640 301.290 286.240 ;
    END
  END A[25]
  PIN A[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 308.010 80.870 312.010 ;
    END
  END A[26]
  PIN A[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END A[27]
  PIN A[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END A[28]
  PIN A[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 119.040 301.290 119.640 ;
    END
  END A[29]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END A[2]
  PIN A[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 170.040 301.290 170.640 ;
    END
  END A[30]
  PIN A[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 91.840 301.290 92.440 ;
    END
  END A[31]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 234.640 301.290 235.240 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 40.840 301.290 41.440 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 272.040 301.290 272.640 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 308.010 190.350 312.010 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 308.010 142.050 312.010 ;
    END
  END B[0]
  PIN B[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END B[10]
  PIN B[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 308.010 251.530 312.010 ;
    END
  END B[11]
  PIN B[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END B[12]
  PIN B[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 0.040 301.290 0.640 ;
    END
  END B[13]
  PIN B[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END B[14]
  PIN B[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 308.010 129.170 312.010 ;
    END
  END B[15]
  PIN B[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 308.010 167.810 312.010 ;
    END
  END B[16]
  PIN B[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 308.010 264.410 312.010 ;
    END
  END B[17]
  PIN B[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END B[18]
  PIN B[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 221.040 301.290 221.640 ;
    END
  END B[19]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END B[1]
  PIN B[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 308.010 180.690 312.010 ;
    END
  END B[20]
  PIN B[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END B[21]
  PIN B[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 54.440 301.290 55.040 ;
    END
  END B[22]
  PIN B[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 156.440 301.290 157.040 ;
    END
  END B[23]
  PIN B[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END B[24]
  PIN B[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END B[25]
  PIN B[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END B[26]
  PIN B[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END B[27]
  PIN B[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END B[28]
  PIN B[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 308.010 32.570 312.010 ;
    END
  END B[29]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END B[2]
  PIN B[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END B[30]
  PIN B[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END B[31]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 129.240 301.290 129.840 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 64.640 301.290 65.240 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 13.640 301.290 14.240 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 308.010 45.450 312.010 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 105.440 301.290 106.040 ;
    END
  END B[9]
  PIN F[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END F[0]
  PIN F[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END F[10]
  PIN F[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 207.440 301.290 208.040 ;
    END
  END F[11]
  PIN F[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 308.010 58.330 312.010 ;
    END
  END F[12]
  PIN F[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END F[13]
  PIN F[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END F[14]
  PIN F[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END F[15]
  PIN F[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END F[16]
  PIN F[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END F[17]
  PIN F[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 308.010 154.930 312.010 ;
    END
  END F[18]
  PIN F[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END F[19]
  PIN F[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 308.010 6.810 312.010 ;
    END
  END F[1]
  PIN F[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END F[20]
  PIN F[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END F[21]
  PIN F[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 308.010 277.290 312.010 ;
    END
  END F[22]
  PIN F[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 308.010 216.110 312.010 ;
    END
  END F[23]
  PIN F[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END F[24]
  PIN F[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 308.010 299.830 312.010 ;
    END
  END F[25]
  PIN F[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 27.240 301.290 27.840 ;
    END
  END F[26]
  PIN F[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END F[27]
  PIN F[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END F[28]
  PIN F[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END F[29]
  PIN F[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END F[2]
  PIN F[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END F[30]
  PIN F[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 183.640 301.290 184.240 ;
    END
  END F[31]
  PIN F[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END F[3]
  PIN F[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 308.010 241.870 312.010 ;
    END
  END F[4]
  PIN F[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 308.010 228.990 312.010 ;
    END
  END F[5]
  PIN F[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 308.010 19.690 312.010 ;
    END
  END F[6]
  PIN F[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 308.010 67.990 312.010 ;
    END
  END F[7]
  PIN F[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END F[8]
  PIN F[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END F[9]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 295.320 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 295.320 257.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 299.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 299.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 295.320 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 295.320 181.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 299.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 299.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 297.290 142.840 301.290 143.440 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 295.320 299.285 ;
      LAYER met1 ;
        RECT 0.070 5.820 299.850 299.840 ;
      LAYER met2 ;
        RECT 0.100 307.730 6.250 309.925 ;
        RECT 7.090 307.730 19.130 309.925 ;
        RECT 19.970 307.730 32.010 309.925 ;
        RECT 32.850 307.730 44.890 309.925 ;
        RECT 45.730 307.730 57.770 309.925 ;
        RECT 58.610 307.730 67.430 309.925 ;
        RECT 68.270 307.730 80.310 309.925 ;
        RECT 81.150 307.730 93.190 309.925 ;
        RECT 94.030 307.730 106.070 309.925 ;
        RECT 106.910 307.730 118.950 309.925 ;
        RECT 119.790 307.730 128.610 309.925 ;
        RECT 129.450 307.730 141.490 309.925 ;
        RECT 142.330 307.730 154.370 309.925 ;
        RECT 155.210 307.730 167.250 309.925 ;
        RECT 168.090 307.730 180.130 309.925 ;
        RECT 180.970 307.730 189.790 309.925 ;
        RECT 190.630 307.730 202.670 309.925 ;
        RECT 203.510 307.730 215.550 309.925 ;
        RECT 216.390 307.730 228.430 309.925 ;
        RECT 229.270 307.730 241.310 309.925 ;
        RECT 242.150 307.730 250.970 309.925 ;
        RECT 251.810 307.730 263.850 309.925 ;
        RECT 264.690 307.730 276.730 309.925 ;
        RECT 277.570 307.730 289.610 309.925 ;
        RECT 290.450 307.730 299.270 309.925 ;
        RECT 0.100 4.280 299.820 307.730 ;
        RECT 0.650 0.155 9.470 4.280 ;
        RECT 10.310 0.155 22.350 4.280 ;
        RECT 23.190 0.155 35.230 4.280 ;
        RECT 36.070 0.155 48.110 4.280 ;
        RECT 48.950 0.155 57.770 4.280 ;
        RECT 58.610 0.155 70.650 4.280 ;
        RECT 71.490 0.155 83.530 4.280 ;
        RECT 84.370 0.155 96.410 4.280 ;
        RECT 97.250 0.155 109.290 4.280 ;
        RECT 110.130 0.155 118.950 4.280 ;
        RECT 119.790 0.155 131.830 4.280 ;
        RECT 132.670 0.155 144.710 4.280 ;
        RECT 145.550 0.155 157.590 4.280 ;
        RECT 158.430 0.155 170.470 4.280 ;
        RECT 171.310 0.155 180.130 4.280 ;
        RECT 180.970 0.155 193.010 4.280 ;
        RECT 193.850 0.155 205.890 4.280 ;
        RECT 206.730 0.155 218.770 4.280 ;
        RECT 219.610 0.155 231.650 4.280 ;
        RECT 232.490 0.155 241.310 4.280 ;
        RECT 242.150 0.155 254.190 4.280 ;
        RECT 255.030 0.155 267.070 4.280 ;
        RECT 267.910 0.155 279.950 4.280 ;
        RECT 280.790 0.155 292.830 4.280 ;
        RECT 293.670 0.155 299.820 4.280 ;
      LAYER met3 ;
        RECT 4.400 309.040 297.290 309.905 ;
        RECT 4.000 300.240 297.290 309.040 ;
        RECT 4.000 298.840 296.890 300.240 ;
        RECT 4.000 296.840 297.290 298.840 ;
        RECT 4.400 295.440 297.290 296.840 ;
        RECT 4.000 286.640 297.290 295.440 ;
        RECT 4.000 285.240 296.890 286.640 ;
        RECT 4.000 283.240 297.290 285.240 ;
        RECT 4.400 281.840 297.290 283.240 ;
        RECT 4.000 273.040 297.290 281.840 ;
        RECT 4.000 271.640 296.890 273.040 ;
        RECT 4.000 269.640 297.290 271.640 ;
        RECT 4.400 268.240 297.290 269.640 ;
        RECT 4.000 259.440 297.290 268.240 ;
        RECT 4.000 258.040 296.890 259.440 ;
        RECT 4.000 256.040 297.290 258.040 ;
        RECT 4.400 254.640 297.290 256.040 ;
        RECT 4.000 249.240 297.290 254.640 ;
        RECT 4.000 247.840 296.890 249.240 ;
        RECT 4.000 245.840 297.290 247.840 ;
        RECT 4.400 244.440 297.290 245.840 ;
        RECT 4.000 235.640 297.290 244.440 ;
        RECT 4.000 234.240 296.890 235.640 ;
        RECT 4.000 232.240 297.290 234.240 ;
        RECT 4.400 230.840 297.290 232.240 ;
        RECT 4.000 222.040 297.290 230.840 ;
        RECT 4.000 220.640 296.890 222.040 ;
        RECT 4.000 218.640 297.290 220.640 ;
        RECT 4.400 217.240 297.290 218.640 ;
        RECT 4.000 208.440 297.290 217.240 ;
        RECT 4.000 207.040 296.890 208.440 ;
        RECT 4.000 205.040 297.290 207.040 ;
        RECT 4.400 203.640 297.290 205.040 ;
        RECT 4.000 194.840 297.290 203.640 ;
        RECT 4.000 193.440 296.890 194.840 ;
        RECT 4.000 191.440 297.290 193.440 ;
        RECT 4.400 190.040 297.290 191.440 ;
        RECT 4.000 184.640 297.290 190.040 ;
        RECT 4.000 183.240 296.890 184.640 ;
        RECT 4.000 181.240 297.290 183.240 ;
        RECT 4.400 179.840 297.290 181.240 ;
        RECT 4.000 171.040 297.290 179.840 ;
        RECT 4.000 169.640 296.890 171.040 ;
        RECT 4.000 167.640 297.290 169.640 ;
        RECT 4.400 166.240 297.290 167.640 ;
        RECT 4.000 157.440 297.290 166.240 ;
        RECT 4.000 156.040 296.890 157.440 ;
        RECT 4.000 154.040 297.290 156.040 ;
        RECT 4.400 152.640 297.290 154.040 ;
        RECT 4.000 143.840 297.290 152.640 ;
        RECT 4.000 142.440 296.890 143.840 ;
        RECT 4.000 140.440 297.290 142.440 ;
        RECT 4.400 139.040 297.290 140.440 ;
        RECT 4.000 130.240 297.290 139.040 ;
        RECT 4.000 128.840 296.890 130.240 ;
        RECT 4.000 126.840 297.290 128.840 ;
        RECT 4.400 125.440 297.290 126.840 ;
        RECT 4.000 120.040 297.290 125.440 ;
        RECT 4.000 118.640 296.890 120.040 ;
        RECT 4.000 116.640 297.290 118.640 ;
        RECT 4.400 115.240 297.290 116.640 ;
        RECT 4.000 106.440 297.290 115.240 ;
        RECT 4.000 105.040 296.890 106.440 ;
        RECT 4.000 103.040 297.290 105.040 ;
        RECT 4.400 101.640 297.290 103.040 ;
        RECT 4.000 92.840 297.290 101.640 ;
        RECT 4.000 91.440 296.890 92.840 ;
        RECT 4.000 89.440 297.290 91.440 ;
        RECT 4.400 88.040 297.290 89.440 ;
        RECT 4.000 79.240 297.290 88.040 ;
        RECT 4.000 77.840 296.890 79.240 ;
        RECT 4.000 75.840 297.290 77.840 ;
        RECT 4.400 74.440 297.290 75.840 ;
        RECT 4.000 65.640 297.290 74.440 ;
        RECT 4.000 64.240 296.890 65.640 ;
        RECT 4.000 62.240 297.290 64.240 ;
        RECT 4.400 60.840 297.290 62.240 ;
        RECT 4.000 55.440 297.290 60.840 ;
        RECT 4.000 54.040 296.890 55.440 ;
        RECT 4.000 52.040 297.290 54.040 ;
        RECT 4.400 50.640 297.290 52.040 ;
        RECT 4.000 41.840 297.290 50.640 ;
        RECT 4.000 40.440 296.890 41.840 ;
        RECT 4.000 38.440 297.290 40.440 ;
        RECT 4.400 37.040 297.290 38.440 ;
        RECT 4.000 28.240 297.290 37.040 ;
        RECT 4.000 26.840 296.890 28.240 ;
        RECT 4.000 24.840 297.290 26.840 ;
        RECT 4.400 23.440 297.290 24.840 ;
        RECT 4.000 14.640 297.290 23.440 ;
        RECT 4.000 13.240 296.890 14.640 ;
        RECT 4.000 11.240 297.290 13.240 ;
        RECT 4.400 9.840 297.290 11.240 ;
        RECT 4.000 1.040 297.290 9.840 ;
        RECT 4.000 0.175 296.890 1.040 ;
      LAYER met4 ;
        RECT 9.495 11.055 20.640 290.185 ;
        RECT 23.040 11.055 97.440 290.185 ;
        RECT 99.840 11.055 174.240 290.185 ;
        RECT 176.640 11.055 251.040 290.185 ;
        RECT 253.440 11.055 275.705 290.185 ;
      LAYER met5 ;
        RECT 75.100 34.900 155.820 53.500 ;
  END
END MULTI_32bit
END LIBRARY

